module uart2

#define	uart2__any()	U2STAbits.URXDA