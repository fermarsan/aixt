module pwm

