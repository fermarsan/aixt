// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fabián A. Rojas Acosta, Alberto Pinzón Valero and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Pin management functions (LQFP32 MiniEVB Nano - LGT8F328P port)
module pin

// in macro defines the pin input mode
#define input  INPUT
#define input_pullup  INPUT_PULLUP

// out macro defines the pin output mode
#define output  OUTPUT

