module uart

fn C.read() u8