// Author: Fernando M. Santa
// Date: 2024
//
// ## Description
// ADC functions
module adc


// adc channels
pub const ch0 = 36
// pub const ch1 = xx
// pub const ch2 = xx
pub const ch3 = 39
pub const ch4 = 32
pub const ch5 = 33
pub const ch6 = 34
pub const ch7 = 35
pub const ch8 = 25