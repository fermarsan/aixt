module pic16f88x

pub const description = 'API for the PIC16F88x family devices'
