module uart

#define	uart.any()	U1STAbits.URXDA