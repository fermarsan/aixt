// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2023-2024
// License: MIT
//
// Description: This is a module to emulate digital pines in console.
#include <stdio.h>
#include <stdlib.h>

__global (
    pins__ = [0, 0, 0, 0, 0, 0, 0, 0]   // virtual pin array
    input__ = 0
)

// pin_update prints the pins table in the command line
fn pin_update() {
    system("clear")
    printf(" Aixt virtual pins     [#] = ON   [ ] = OFF\n")
    printf(" _____ _____ _____ _____ _____ _____ _____ _____\n")
    printf("|  a  |  b  |  c  |  d  |  w  |  x  |  y  |  z  |\n")
    for i__ := 0; i__<=7; i__++ {
        if pins__[i__] == 0 {
            printf("| [ ] ")
        } else {
            printf("| [#] ")
        }
    }
    printf("|\n'-----'-----'-----'-----'-----'-----'-----'-----'\n")
}

// fn pin_name(pin int) &char {
//     switch (pin) {
//     case a:  return "a";
//     case b:  return "b";
//     case c:  return "c";
//     case d:  return "d";
//     case w:  return "w";
//     case x:  return "x";
//     case y:  return "y";
//     case z:  return "z";    
//     default: return "ERROR";
//     }
// } 

fn pin_high(pin int) {   
   pins__[pin] = 1
    pin_update()
}

fn pin_low(pin int) {   
   pins__[pin] = 0
    pin_update()
}

fn pin_write(pin int, val int) {  
   pins__[pin] = val
    pin_update()
}

fn pin_read(pin  int) int {
    system("clear")
    printf(" Aixt virtual pins     Input %s : ", pin_name(pin))
    scanf("%d", &input__)
    pin_write(pin, input__)
    return input__
}