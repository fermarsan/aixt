// Project name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: delay functions for XC8 compiler

module time

fn C.__delay_ms(tms u16)
fn C.__delay_us(tus u16)