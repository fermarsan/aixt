module uart
#define uart__println_1(MESSAGE)		Serial.println(MESSAGE)

