// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git
// File Name: setup.c.v
// Author: Fernando Martinez Santa - Arley Junco - Luis Quevedo 
// Date: 2024
// License : MIT

module pin 

#define pin__setup(PIN_NAME, MODE)        pinMode(PIN_NAME, MODE)