// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: PWM functions (Explorer16-PIC24 port)
module pwm

#define		pwm__out_1		1
#define		pwm__out_2		2
#define		pwm__out_1_2	3
