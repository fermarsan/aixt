module pic16f6xx_18p

pub const description = 'API for the PIC16f6xx_18p family devices'
