module pic18

pub const description = 'API for the PIC18 family devices'
