// File: https://github.com/fermarsan/aixt/blob/main/
// Author: Fernando M. Santa - Daniel Polo - Edwin Barrera - Javier Leon - Camilo Lucas
// Date: 2022-2025
//
// // ## Description
// time functions (CY8CKIT-145-40XX)

module time


fn C.CyDelay(tms any)
fn C.CyDelayUs(tus any)
