// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: usb_uart module (Arduino Nano - ATmega328P port)
module usb_uart


