module main

#include "CH57x_common.h"
#define true 1

