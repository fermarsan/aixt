// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: pin.c.v
// Author: Fernando Martínez Santa - Johann Escobar Guzmán - Daniel Andrés Vásquez Gómez
// Date: 2023-2024
// License: MIT
//
// // Description: PIN functions (W801)
//              (PC port) 

module pin
#define pwm.pin[PIN_NAME]  pwm_pin[PIN_NAME]