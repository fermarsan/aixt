module main

#include "CH82x_common.h"
#define true 1
