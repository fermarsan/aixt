// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: ADC functions
module adc

fn C.analogReadResolution(res any)

// adc channels
pub const ch0 = A0
pub const ch1 = A1
pub const ch2 = A2
pub const ch3 = A3
pub const ch4 = A4
pub const ch5 = A5
pub const ch6 = A6
pub const ch7 = A7
