module pwm

fn init(){

}