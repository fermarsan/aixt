// Author: Jan Carlo Peñuela Jurado and Fernando M. Santa
// Date: 2024
//
// ## Description
// uart
//              (PIC18F452)
module uart

#include <xc.h>
