// Project Name : Aixt: http://github.com/fermansan/aixt.git
// Authors:
//  - Arley Junco
//  - Luis Quevedo
//  - Fernando M. Santa
//
// _Date:_ 2024
// License : MIT

module pwm

// TODO: PWM channels defining