// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa & Cristian Garzón
// Date: 2023 - 2024
// Description: TIME functions (WCH-CH573F)

module time

#include "CH57x_common.h"

fn init() {

}