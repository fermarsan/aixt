module my_mod

// add (integer)
pub fn add(x int, y int) int {
	return x + y
}