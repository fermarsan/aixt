// Project name: Aixt https://github.com/fermarsan/aixt.git
// Authors: Fernando M. Santa
// Date: 2025
// License: MIT
//
// Description: Builtin LEDs
module leds



