// _File:_ https://github.com/fermarsan/aixt/blob/main/
// Authors:
//	 - Julian Camilo Guzmán Zambrano
//	 - Juan Pablo Gonzalez Penagos
//	 - Fernando M. Santa
//
// _Date:_ 2022-2024
//
// // ## Description
// PWM functions (Blue Pill_STM32F103C)
//              (PC port)

module pwm

@[inline]
pub fn write(PIN_NAME, MODE) {
	C.pwmWrite(PIN_NAME, MODE)
}

@[inline]
pub fn map(MODE, VALUE,VALUE1,VALUE2,VALUE3) {
	C.map(MODE, VALUE,VALUE1,VALUE2,VALUE3)
}
