// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: ADC functions
module adc

fn C.analogReadResolution(res any)	

// adc channels
pub const ch0 = 36
// pub const ch1 = xx
// pub const ch2 = xx
pub const ch3 = 39
pub const ch4 = 32
pub const ch5 = 33
pub const ch6 = 34
pub const ch7 = 35
pub const ch8 = 25