// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fabián A. Rojas Acosta, Alberto Pinzón Valero and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: Pin management functions (LQFP32 MiniEVB Nano - LGT8F328P port)
module pin

// in macro defines the pin input mode
#define pin__input  INPUT
#define pin__input_pullup  INPUT_PULLUP

// out macro defines the pin output mode
#define pin__output  OUTPUT

fn init() { //  init function call setup or initialization code

}