// Project Name : Aixt: http://github.com/fermansan/aixt.git
// Authors:
//  - Arley Junco
//  - Luis Quevedo
//  - Fernando M. Santa
// Date: 2024
// License : MIT

module time

#define time.sleep(S)   delay(S*1000)

#define time.sleep_ms(MS)  delay(MS)

#define time.sleep_us(US)   delayMicroseconds(US)