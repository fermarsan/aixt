module pin

#define pin.low(PIN_NAME)		digitalWrite(PIN_NAME, LOW)
