// Project name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2025
// License: MIT
//
// Description: Pin management functions for 16F family
module pin

#include "low_fast.c"

fn C.LOW_FAST(port_name u8, pin_number u8)

// low_fast puts a logic 1 to a pin faster than the low function
@[as_macro]
pub fn low_fast(port_name u8, pin_number u8) {
	C.LOW_FAST(port_name, pin_number)
}
