// _File:_ https://github.com/fermarsan/aixt/blob/main/
//
// _Authors:_ Fernando M. Santa
//
// _Date:_ 2025
//
// ## Description
// Builtin definitions PIC12F6xx

module main

#include <xc.h>
#include <stdint.h>
#include <stdbool.h>

#include "builtin.c"
