// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Cristian Garzón
// Date: 2023 - 2024
// Description: UART functions (WCH-CH582F)

module uart 

#define uart.println(MSG)		uart.print(MSG);  uart.write('\n');  uart.write('\r')