// module importing

import time { sleep }
import machine

a := 0

for {
	sleep(1)
	a++
}