// Author: Fernando M. Santa
// Date: 2022-2025
//
// ## Description
// Builtin definitions (STM32F411Core port)
module main
