// Author: Cristian Garzón
// Date: 2023 - 2024
// ## Description
// UART functions (WCH-CH582F)

module uart

fn C.read() u8
