module xc8

pub const description = 'Workspace for the xc8 compiler modules'
