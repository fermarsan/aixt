// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// File Name: pin.c.v
// Author: Andrés Felipe Fajardo Duarte and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: PIN management functions  (PIC18F2550 port)

module pin

#include <xc.h>

#define pin__output  0   // pin mode (direction)
#define pin__input   1

fn init() {

}