module uno

pub const description = 'Arduino Uno target API'
