// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2022-2024
//
// ## Description
// Builtin definitions (Exp16-PIC24 port)
module main

#include <xc.h>
#include <stdint.h>
#include <stdbool.h>

#include "builtin.c"




// fn C.init()