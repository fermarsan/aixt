module pwm

fn init() {

}