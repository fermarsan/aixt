// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2022-2024
// License: MIT
module time

// sleep_us is a delay function in microseconds for the Aixt Exp16-PIC24 port. 
#define time.sleep_us(TIME)    __delay_us(TIME)