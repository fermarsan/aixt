module time

#define time.sleep_us(TIME)	delayMicroseconds(TIME)
