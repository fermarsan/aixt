// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: dutymin.c.v
// Author: Fernando M. Santa - Johann Escobar Guzmán - Daniel Andrés Vásquez Gómez
// Date: 2023-2024
// License: MIT
//
// // Description: DUTY_MIN functions (W801)
//              (PC port) 

module pin

#define DUTY__MIN  DUTY_MIN