module PIC12

pub const description = 'Workspace for the PIC12 family devices'
