// Project name: Aixt, https://github.com/fermarsan/aixt.git
//
// _Author:_ Fernando M. Santa
//
// _Date:_ 2024
// License: MIT

// module uart

// any function gets the number of bytes (characters) available for reading
// @[as_macro]
// pub fn any() int {
// 	return C.SERIAL_AVAILABLE()
// }
