// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git

// Author: Farith Ochoa León, Delipe Cardozo and Fernando M. Santa 
// License : MIT

module pin 

#define pin.setup(PIN_NAME, MODE) 	 	 pinMode(PIN_NAME, MODE)