// Author: Fernando M. Santa
// Date: 2024


// module uart

// any function gets the number of bytes (characters) available for reading
// @[as_macro]
// pub fn any() int {
// 	return C.SERIAL_AVAILABLE()
// }
