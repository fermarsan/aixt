// _File:_ https://github.com/fermarsan/aixt/blob/main/
//
// _Author:_ Fernando M. Santa
//
// _Date:_ 2022-2025
//
// ## Description
// Builtin definitions (XIAO-SAMD21 port)
module main
