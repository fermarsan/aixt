module pin

#define pin.high(PIN_NAME)		digitalWrite(PIN_NAME, HIGH)
