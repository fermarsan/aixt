module adc