// Author: Fernando M. Santa
// Date: 2024-2025
//
// ## Description
// ADC functions
module adc

// adc channels
pub const ch0 = 26
pub const ch1 = 27
pub const ch2 = 28