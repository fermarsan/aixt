module pin

#define pin__high(PIN_NAME)		digitalWrite(PIN_NAME, HIGH)
fn_init(){

}