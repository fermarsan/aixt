module xc16

pub const description = 'API for the xc16 compiler modules'
