module pin

#define pin__write(PIN_NAME, VALUE)		digitalWrite(PIN_NAME, VALUE)