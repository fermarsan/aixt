// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2025
//
// ## Description
// Random numbers functions
module random

#include "random.c"

fn C.RANDOMINRANGE(min int, max int) int
fn C.random(max int) int
fn C.randomSeed(s u32)