module uart

#define uart__ready_1()		Serial1.available()