// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fabián A. Rojas Acosta, Alberto Pinzón Valero and Fernando M. Santa
// Date: 2024
// License: MIT
module time

//Pauses the program for the amount of time (in microseconds) specified by the parameter
#define time.sleep_us(TUS)  delayMicroseconds(TUS)