// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: ADC functions Arduinio Uno
module adc_fn

// ADC pin names
@[as_macro] pub const ch0 = 54
@[as_macro] pub const ch1 = 55
@[as_macro] pub const ch2 = 56
@[as_macro] pub const ch3 = 57
@[as_macro] pub const ch4 = 58
@[as_macro] pub const ch5 = 59
@[as_macro] pub const ch6 = 60
@[as_macro] pub const ch7 = 61
@[as_macro] pub const ch8 = 62
@[as_macro] pub const ch9 = 63
@[as_macro] pub const ch10 = 64
@[as_macro] pub const ch11 = 65
@[as_macro] pub const ch12 = 66
@[as_macro] pub const ch13 = 67
@[as_macro] pub const ch14 = 68
@[as_macro] pub const ch15 = 69
