// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// File Name: uart setup.c.v
// Author: Luis Alfredo Pinto Medina and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Pin management functions
//              (PIC16F886 port)

module uart

fn C.setup(baudrate u32)