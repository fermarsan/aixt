module core

pub const description = 'Arduino core API'
