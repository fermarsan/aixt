module xc8

pub const description = 'API for the xc8 compiler modules'
