// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: builtin.c
// Author: Fernando Martínez Santa - Julian Camilo Guzmán Zambrano - Juan Pablo Gonzalez Penagos
// Date: 2022-2023
// License: MIT
//
// Description: Builtin definitions
//              (PC port) 
module main

enum __pin_names {    // enumerated type for the pin names
 
    rx=PA9
    tx=PA10
    p1=PA0
    p2=PA1
    p3=PA2
    p4=PA3
    p5=PA4
    p6=PA5
    p7=PA6
    p8=PA7
    p9=PA8
    p10=PA13
    p11=PA14
    p12=PA15
    p13=PB0
    p14=PB1
    p15=PB2
    p16=PB3
    p17=PB4
    p18=PB5
    p19=PB6
    p20=PB7
    p21=PB8
    p22=PB9
    p23=PB10
    p24=PB11
    p25=PB12
    p26=PB13
    p27=PB14
    p28=PB15

recibe_dato
dato
envia_dato
}



fn init() {

}
