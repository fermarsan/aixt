// Project name: Aixt, https://github.com/fermarsan/aixt.git
//
// _Author:_ Jan Carlo Peñuela Jurado and Fernando M. Santa
//
// _Date:_ 2024
//
// ## Description
// PWM WRITE
//              (PIC18F452)
module pwm
fn write(duty int)    
    { 
        pwm := ((duty - 0) * (50 - 0) / (1023 - 0) + 0) /* Calculando el ciclo de trabajo */ 
        CCPR1L = pwm >> 2 /* Almacena el valor del PWM */ 
    }