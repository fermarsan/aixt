// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Pin management functions Arduino devices
module pin

// pin names
// @[as_macro] pub const pa0   = 0    
@[as_macro] pub const a1   = u8(C.PA1) 
@[as_macro] pub const a2   = u8(C.PA2) 
@[as_macro] pub const a3   = u8(C.PA3) 
@[as_macro] pub const a4   = u8(C.PA4) 
@[as_macro] pub const a5   = u8(C.PA5) 
@[as_macro] pub const a6   = u8(C.PA6) 
@[as_macro] pub const a7   = u8(C.PA7) 
@[as_macro] pub const a8   = u8(C.PA8) 
@[as_macro] pub const a9   = u8(C.PA9) 
@[as_macro] pub const a10  = u8(C.PA10)
@[as_macro] pub const a11  = u8(C.PA11)
@[as_macro] pub const a12  = u8(C.PA12)
@[as_macro] pub const a13  = u8(C.PA13)
@[as_macro] pub const a14  = u8(C.PA14)
@[as_macro] pub const a15  = u8(C.PA15)

@[as_macro] pub const b0   = u8(C.PB0)   
@[as_macro] pub const b1   = u8(C.PB1) 
@[as_macro] pub const b2   = u8(C.PB2) 
@[as_macro] pub const b3   = u8(C.PB3) 
@[as_macro] pub const b4   = u8(C.PB4) 
@[as_macro] pub const b5   = u8(C.PB5) 
@[as_macro] pub const b6   = u8(C.PB6) 
@[as_macro] pub const b7   = u8(C.PB7) 
@[as_macro] pub const b8   = u8(C.PB8) 
@[as_macro] pub const b9   = u8(C.PB9) 
@[as_macro] pub const b10  = u8(C.PB10)
@[as_macro] pub const b11  = u8(C.PB11)
@[as_macro] pub const b12  = u8(C.PB12)
@[as_macro] pub const b13  = u8(C.PB13)
@[as_macro] pub const b14  = u8(C.PB14)
@[as_macro] pub const b15  = u8(C.PB15)
@[as_macro] pub const b16  = u8(C.PB16)
@[as_macro] pub const b17  = u8(C.PB17)
@[as_macro] pub const b18  = u8(C.PB18)
@[as_macro] pub const b19  = u8(C.PB19)
@[as_macro] pub const b20  = u8(C.PB20)
@[as_macro] pub const b21  = u8(C.PB21)
@[as_macro] pub const b22  = u8(C.PB22)
@[as_macro] pub const b23  = u8(C.PB23)
@[as_macro] pub const b24  = u8(C.PB24)
@[as_macro] pub const b25  = u8(C.PB25)
@[as_macro] pub const b26  = u8(C.PB26)
@[as_macro] pub const b27  = u8(C.PB27)
