module adc

#define adc__write(PIN_NAME)   analogWrite(PIN_NAME)