module PIC24_dsPIC33

pub const description = 'Workspace for the PIC24_dsPIC33 family devices'
