module arduino

pub const description = 'Arduino targets API'
