module main

import my_mod.my_sub

fn main() {
	my_sub.add(3,4)
	my_sub.sub(23,21)
}