// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git

// Author: Fernando M. Santa - Arley Junco - Luis Quevedo 
// Date: 2024
// License : MIT


module adc 

#define adc__read(PIN_NAME)    analogRead(PIN_NAME)