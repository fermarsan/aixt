// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: PWM functions (Explorer16-PIC24 port)
module pwm

#define		pwm.out_1		1
#define		pwm.out_2		2
#define		pwm.out_1_2	3
