// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Pin management functions Arduino devices
module pin

// pin names
// pub const pa0   = 0    
pub const a1   = C.PA1 
pub const a2   = C.PA2 
pub const a3   = C.PA3 
pub const a4   = C.PA4 
pub const a5   = C.PA5 
pub const a6   = C.PA6 
pub const a7   = C.PA7 
pub const a8   = C.PA8 
pub const a9   = C.PA9 
pub const a10  = C.PA10
pub const a11  = C.PA11
pub const a12  = C.PA12
pub const a13  = C.PA13
pub const a14  = C.PA14
pub const a15  = C.PA15

pub const b0   = C.PB0   
pub const b1   = C.PB1 
pub const b2   = C.PB2 
pub const b3   = C.PB3 
pub const b4   = C.PB4 
pub const b5   = C.PB5 
pub const b6   = C.PB6 
pub const b7   = C.PB7 
pub const b8   = C.PB8 
pub const b9   = C.PB9 
pub const b10  = C.PB10
pub const b11  = C.PB11
pub const b12  = C.PB12
pub const b13  = C.PB13
pub const b14  = C.PB14
pub const b15  = C.PB15
pub const b16  = C.PB16
pub const b17  = C.PB17
pub const b18  = C.PB18
pub const b19  = C.PB19
pub const b20  = C.PB20
pub const b21  = C.PB21
pub const b22  = C.PB22
pub const b23  = C.PB23
pub const b24  = C.PB24
pub const b25  = C.PB25
pub const b26  = C.PB26
pub const b27  = C.PB27

// pin modes
pub const input		= 0
pub const output	= 1
pub const in_pullup = 2
