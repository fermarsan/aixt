// Author: Fernando M. Santa
// Date: 2024-2025
//
// ## Description
// UART module (Arduino Nano - ATmega328P port)
module uart

// NOTE: this is the USB-UART, you could import it like:
//		`import uart as usb_uart`

