// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fabián A. Rojas Acosta, Alberto Pinzón Valero and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: ADC functions (LQFP32 MiniEVB Nano - LGT8F328P port)
module adc

// define analog pins
@[as_macro] pub const a0 =  A0  
@[as_macro] pub const a1 =  A1
@[as_macro] pub const a2 =  A2
@[as_macro] pub const a3 =  A3
@[as_macro] pub const a4 =  A4
@[as_macro] pub const a5 =  A5
@[as_macro] pub const a6 =  A6
@[as_macro] pub const a7 =  A7
@[as_macro] pub const a10 =  A10