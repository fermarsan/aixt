module cypress

pub const description = 'Cypress targets API'
