// Author: Cristian Garzón
// Date: 2023 - 2024
// ## Description
// UART functions (WCH-CH573F)

module uart

fn C.setup(baud_rate u32)
