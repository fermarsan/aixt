module uart
#define uart.write(VALUE)    Serial.write(VALUE)