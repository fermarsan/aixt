// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git
// File Name: sleep.c.v
// Author: Fernando Martinez Santa - Arley Junco - Luis Quevedo 
// Date: 2024
// License : MIT

module time

#define time__sleep(S)   delay(S*1000)
