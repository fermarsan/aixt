module equivalents

pub const dict := {
	'x':	'X'
	'y':	'YY'
	'z':	'ZZZ'
}