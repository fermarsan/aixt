// Author: Fernando M. Santa
// Date: 2024
//
// ## Description
// PWM functions (Exp16-PIC24 port)
module pwm

#define		pwm.out_1		1
#define		pwm.out_2		2
#define		pwm.out_1_2	3
