// Project name: Aixt, https://github.com/fermarsan/aixt.git
//
// _Author:_ Fernando M. Santa
//
// _Date:_ 2024
//
// ## Description
// PWM functions (Arduino Nano - ATmega328P port)
module pwm

fn C.analogwrite(id u8, value u8)