// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: write.c.v
// Author: Fernando Martínez Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: WRITE functions (Ai_Thinker_Ai-WB2-32S-Kit)
//              (PC port) 

module adc

#define adc__write(PIN_NAME)   analogWrite(PIN_NAME)