
module pin

#define pin__setup(PIN_NAME, MODE)    pinMode(PIN_NAME, MODE)