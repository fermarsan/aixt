// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// File Name: read.c.v
// Author: Jan Carlo Peñuela Jurado and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: read UART
//              (PIC18F452)
module uart

fn read() rune{
  return RCREG  
}