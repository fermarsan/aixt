// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fabián A. Rojas Acosta, Alberto Pinzón Valero and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: ADC functions (Arduino Nano - ATmega328P port)
module adc

fn init() { //  init function call setup or initialization code

}