// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2022-2024
// License: MIT
module time

#include <unistd.h>

// sleep is a delay function in seconds for the Aixt PC port. 
#define time__sleep(TIME)		sleep(TIME)