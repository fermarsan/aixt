// Project Name: Aixt project, https://gitlab.com/fermarsan/aixt-project.git
// File Name: pin.c.v
// Author: Jan Carlo Peñuela Jurado and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: Pin management functions (PIC18F452)
module pin

#include <xc.h>

#define pin__output 0   // pin mode (direction)
#define pin__input  1

fn init() {
    
}