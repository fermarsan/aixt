// Project name: Aixt, https://github.com/fermarsan/aixt.git
//
// _Author:_ Fabián A. Rojas Acosta, Alberto Pinzón Valero and Fernando M. Santa
//
// _Date:_ 2024
//
// ## Description
// PWM functions (LQFP32 MiniEVB Nano - LGT8F328P port)
module pwm

// TODO: PWM channels defining

