// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fabián A. Rojas Acosta, Alberto Pinzón Valero and Fernando Martínez Santa
// Date: 2024
// License: MIT
module pin

//Write a HIGH or a LOW value to a digital pin
#define pin__write(PIN_NAME, VALUE)  digitalWrite(PIN_NAME, VALUE)  