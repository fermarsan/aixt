// _File:_ https://github.com/fermarsan/aixt/blob/main/
//
// _Author:_ Fernando M. Santa - Daniel Polo - Edwin Barrera - Javier Leon - Camilo Lucas
//
// _Date:_ 2022-2025
//
// // ## Description
// pin functions (CY8CKIT-049-42XX)

module pin

#include "pin.c"


fn C.PIN_WRITE(name any, value any)
fn C.PIN_HIGH(name any)
fn C.PIN_LOW(name any)
fn C.PIN_READ(name any) u8
