// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2022-2024
// License: MIT
//
// Description: Milliseconds delay function
//              (Explorer16-PIC24 port)
module time

#include <libpic30.h>
