// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Cristian Garzón
// Date: 2023 - 2024
// Description: ADC functions (WCH-CH582F)

module adc

#define adc__setup(channel)  ADC_ChannelCfg(channel)

