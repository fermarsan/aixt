// Project Name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Luis Alfredo Pinto Medina and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: Pin-port functions (PIC16F84A port)

module port

#define TRISa	TRISA	// port setup name equivalents
#define TRISb	TRISB

#define PORTa	PORTA	// port in name equivalents
#define PORTb	PORTB

