module uart