// Project Name : Aixt: http://github.com/fermansan/aixt.git
// Author: Fernando M. Santa 
// License : MIT
// Date: 2025
//
// ## Description
// Pin management functions ESP32C3-CORE
module pin

// pin names 
pub const gp0 = 0 
pub const gp1 = 1
pub const gp2 = 2
pub const gp3 = 3
pub const gp4 = 4
pub const gp5 = 5
pub const gp6 = 6
pub const gp7 = 7
pub const gp8 = 8
pub const gp9 = 9
pub const gp10 = 10
pub const gp11 = 11
pub const gp12 = 12
pub const gp13 = 13

pub const gp18 = 18
pub const gp19 = 19