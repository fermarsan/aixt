// Project Name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: External interrupts management functions for 16F family
module ext_irq

#include "ext.c"

@[as_macro] pub const rising =	1
@[as_macro] pub const falling = 0