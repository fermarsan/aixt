// Project name: Aixt, https://github.com/fermarsan/aixt.git
//
// _Author:_ Cristian Garzón
//
// _Date:_ 2023 - 2024
// ## Description
// TIME functions (WCH-CH573F)

module time

#define time.sleep_ms(TIME)    DelayMs(TIME)

