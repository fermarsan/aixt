// Project Name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Luis Alfredo Pinto Medina and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: Pin-port functions (PIC16F8x port)
module port

enum port__names as u8 {
	a = 0
	b =
	c =
	d =
	e = 
}
