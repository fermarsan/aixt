// _File:_ https://github.com/fermarsan/aixt/blob/main/
//
// _Author:_ Cesar Alejandro Roa Acosta and Fernando M. Santa
//
// _Date:_ 2024-2025
//
// ## Description
// Builtin definitions
//              (PIC16F87x)
module main

#include <xc.h>
#include <stdbool.h>
#include <stdint.h>

#include "builtin.c"
