// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git
// File Name: adc.c.v
// Author: Farith Ochoa León, Delipe Cardozo and Fernando Martinez Santa 
// License : MIT

module pwm 

fn init() {

}