// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: time.c.v
// Author: Fernando Martínez Santa - Julian Camilo Guzmán Zambrano - Juan Pablo Gonzalez Penagos
// Date: 2022-2024
// License: MIT
//
// // Description: TIME functions (Blue Pill_STM32F103C)
//              (PC port) 

module time

fn init() {
	
}