// _File:_ https://github.com/fermarsan/aixt/blob/main/
// Authors:
//	- Luis Alfredo Pinto Medina
//	- Fernando M. Santa
//
// _Date:_ 2024
//
// ## Description
// Builtin definitions (PIC16F8x port)

module main

#include <xc.h>
#include <stdint.h>
#include <stdbool.h>

#include "builtin.c"
