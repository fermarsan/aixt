module pin

#define pin__read(PIN_NAME)		digitalRead(PIN_NAME)
