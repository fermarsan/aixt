module rune

// ctype.h
#define     rune__is_upper(...)  isupper(__VA_ARGS__)
#define     rune__is_lower(...)  islower(__VA_ARGS__)
#define     rune__is_alpha(...)  isalpha(__VA_ARGS__)
#define     rune__is_digit(...)  isdigit(__VA_ARGS__)
#define     rune__is_alnum(...)  isalnum(__VA_ARGS__)
#define     rune__is_space(...)  isspace(__VA_ARGS__)
#define     rune__is_cntrl(...)  iscntrl(__VA_ARGS__)
#define     rune__is_print(...)  isprint(__VA_ARGS__)
#define     rune__is_graph(...)  isgraph(__VA_ARGS__)
#define     rune__is_punct(...)  ispunct(__VA_ARGS__)
#define     rune__is_xdigit(...) isxdigit(__VA_ARGS__)
#define     rune__to_upper(...)  toupper(__VA_ARGS__)
#define     rune__to_lower(...)  tolower(__VA_ARGS__)
