module pic16f6xx_14p

pub const description = 'API for the PIC16F6xx_14p family devices'
