// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Pin management XIAO-ESP32-xx
module pin

// pin names
pub const d0   = u8(C.D0)    
pub const d1   = u8(C.D1)
pub const d2   = u8(C.D2)
pub const d3   = u8(C.D3)
pub const d4   = u8(C.D4)
pub const d5   = u8(C.D5)
pub const d6   = u8(C.D6)
pub const d7   = u8(C.D7)
pub const d8   = u8(C.D8)
pub const d9   = u8(C.D9)
pub const d10  = u8(C.D10)
