module my_mod

// sub (integer)
pub fn sub(x int, y int) int {
	return x - y
}