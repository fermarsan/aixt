// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git
// File Name: builtin.c
// Author: Fernando Martinez Santa - Arley Junco - Luis Quevedo 
// Date: 2024
// License : MIT
//
//Description: Builtin definitions
//           (PC port)

module main

//#define led		0

//enum __pin_names {    //enumerated type for the pin names 

// GPIO general propouse input output



//-1      //A4, ADC4
//-2	    //A3, ADC3
//-3      //A2, ADC2
//-4      //A1, ADC1
//-5 	    //AO, ADC0
//0 	 	//D0, A5, ADC5
//1		//D1, A6, ADC6
//2  		//D2, A7, ADC7
//3		//D3
//4		//D4
//5		//D5
//6		//D6
//7		//D7
//8		//D8
//9		//D9  PWM
//10		//D10 PWM SS
//11		//D11 MOSI
//12		//D12 MISO
//13		//D13 CSK
//14		//D14
//15		//D15
//16		//D16
//17 		//D19 
//18		//D20 
//19		//D21 
//20		//D22 
//21		//D23  
//22		//D24  
//23		//D17 
//24		//D18 
//25      //

//}  

fn init () {

}