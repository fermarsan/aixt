module main

fn init{
	
}