// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2025
// License: MIT
//
// Description: lcd module (Arduino Nano - ATmega328P port)
module disp7seg

#include "disp7seg.c"


fn C.DISP7SEG_BEGIN() void
fn C.DISP7SEG_SETVALUE(p1 int) 
fn C.DISP7SEG_SETPRECISION(p1 int) 
fn C.DISP7SEG_SETLEADINGZEROS(p1 bool) 
fn C.DISP7SEG_SETBLANK(p1 bool) 
fn C.DISP7SEG_SETDIGIT(p1 int, p2 int) 
fn C.DISP7SEG_SETDECIMALPOINT(p1 int, p2 bool) 





