// Project Name : Aixt: http://github.com/fermansan/aixt.git
// Author: Farith Ochoa León, Delipe Cardozo and Fernando M. Santa 
// License : MIT
// Date: 2024-2025
//
// ## Description
// ADC functions
module adc2

// ADC pin names
pub const ch0 = 5