module main

#include <bflb_platform.h>
#include <hal_gpio.h>
/* USB STDIO */
#include <usb_stdio.h>
#include "io_def.h"

#define led_b	LED_B_PIN
#define led_g	LED_G_PIN
#define led_r	LED_R_PIN


