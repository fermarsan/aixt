// _File:_ https://github.com/fermarsan/aixt/blob/main/
//
// _Author:_ Fernando M. Santa
//
// _Date:_ 2022-2023
//
// ## Description
// Builtin definitions
//              (PC port)
module main

// builtin LED
const led0 = 25
