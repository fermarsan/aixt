module pwm
fn init(){

}