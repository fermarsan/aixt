module uart

#define	uart.any()		RCIF