module time

#define time.sleep_us(US)    delayMicroseconds(US)