// module importing

import time { sleep }
import uart

a := 0.0

for {
	sleep(1)
	a++
}