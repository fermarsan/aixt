module main

fn init() {

}

