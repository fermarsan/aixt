module timer2

