// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: PWM functions W801
module pwm

pub const ch0_0 = C.PA2
pub const ch0_1 = C.PA10
pub const ch0_2 = C.PB0
pub const ch0_3 = C.PB12
pub const ch0_4 = C.PB19

pub const ch1_0 = C.PA3
pub const ch1_1 = C.PA11
pub const ch1_2 = C.PB1
pub const ch1_3 = C.PB13
pub const ch1_4 = C.PB20

pub const ch2_0 = C.PA0
pub const ch2_1 = C.PA12
pub const ch2_2 = C.PB2
pub const ch2_3 = C.PB14
pub const ch2_4 = C.PB24

pub const ch3_0 = C.PA1
pub const ch3_1 = C.PA13
pub const ch3_2 = C.PB3
pub const ch3_3 = C.PB15
pub const ch3_4 = C.PB25

pub const ch4_0 = C.PA4
pub const ch4_1 = C.PA7
pub const ch4_2 = C.PA14
pub const ch4_3 = C.PB16
pub const ch4_4 = C.PB26