// Project Name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: Builtin definitions

module main

enum __pin_names {    // enumerated type for the pin names
   	gpio11=11
   	gpio14=14
   	gpio17=17
   	gpio3=3
   	gpio4=4
   	gpio5=5
   	gpio7=7
   	gpio16=16
   	gpio12=12
}


