// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: pwm.c.v
// Author: Fernando M. Santa - Julian Camilo Guzmán Zambrano - Juan Pablo Gonzalez Penagos
// Date: 2022-2024
// License: MIT
//
// // Description: PWM functions (Blue-Pill)
//              (PC port) 

module pwm

fn init() {

}