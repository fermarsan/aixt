// Project Name: Aixt project, https://gitlab.com/fermarsan/aixt-project.git
// File Name: time.c.v
// Author: Andrés Felipe Fajardo Duarte and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: TIME delay function
//              (PIC18F2550)

module time

#include <xc.h>