// _File:_ https://github.com/fermarsan/aixt/blob/main/
//
// _Author:_ Fernando M. Santa
//
// _Date:_ 2025
//
// ## Description
// External interrupts management functions for the PIC16F family.
module extb

#include "extb.c"
