// Author: Fernando M. Santa
// Date: 2022-2025
//
// ## Description
// Builtin definitions (XIAO-ESP32-xx port)
module main
