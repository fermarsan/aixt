module mega

pub const description = 'Arduino Mega target API'
