module pin

#define output		OUTPUT
#define input		INPUT
#define in_pullup	INPUT_PULLUP

fn init() {

}