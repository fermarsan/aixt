// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa & Cristian Garzón
// Date: 2023 - 2024

module time

// sleep_us is a delay function in microseconds for the (WCH-CH582F)

#define time__sleep_us(TIME)    DelayUs(TIME)

