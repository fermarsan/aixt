module pin

@[inline]
pub fn setup(pin u8, mode u8) {
	C.gpio_set_mode(pin, mode)
}
