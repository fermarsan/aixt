// Project name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Cesar Alejandro Roa Acosta and Fernando M. Santa
// Date: 2024-2025
// License: MIT
//
// Description: Builtin definitions
//              (PIC16F676)
module main

#include <xc.h>
#include <stdbool.h>
#include <stdint.h>

#include "builtin.C"