// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git

// Author: Farith Ochoa León, Delipe Cardozo and Fernando M. Santa 
// License : MIT

module pin 

#define pin__high(PIN_NAME) 	 	digitalWrite(PIN_NAME, HIGH)