module adc
fn.init(){

}