// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Cristian Garzón
// Date: 2023 - 2024
// Description: UART3 functions (WCH-CH573F)

module uart3

#define uart3__println(MSG)		uart3__print(MSG);  uart3__write('\n');  uart3__write('\r')