// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git
// File Name: builtin.c.v
// Author: Farith Ochoa Leon, Felipe Cardozo and Fernando M. Santa
// Date: 2024
// License : MIT
//
//Description: Builtin definitions (ESP32-C3FH4)
//           

module main

fn init () {

}