module pic24

pub const description = 'API for the PIC24 family devices'
