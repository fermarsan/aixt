module pin

#define pin__write(PIN, VALUE)	gpio_write(PIN, VALUE)