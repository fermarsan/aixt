// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// File Name: uart.c.v
// Author: Cesar Alejandro Roa Acosta and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Uart management functions
//              (PIC16F873A port)

module uart

fn init() {
    
}