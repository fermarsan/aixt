// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2022-2024
// License: MIT
module main

#include <stdbool.h>

// Pin_names is the enumerated type for the pin names
enum Pin_names {
    a = 0   
    b
    c
    d
    w
    x
    y
    z
}

// Channel_names is the enumerated type for the ADC channel names
enum Channel_names {
    ch_0 = 0
    ch_1   
}

// init function call setup or initialization code
fn init() {
    // my_var := 3.45
}