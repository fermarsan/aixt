// Project name: Aixt, https://github.com/fermarsan/aixt.git
//
// _Author:_ Andrés Felipe Fajardo y Fernando M. Santa
//
// _Date:_ 2024
//
// ## Description
// Pin port management functions (PIC18F2550 port)

module port

#include <xc.h>

const output = C.0   // port mode (direction)
const input = C.1


