module uart2

#define	uart2.any()	U2STAbits.URXDA