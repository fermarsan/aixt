// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: builtin.c
// Author: Fernando Martínez Santa - Julian Camilo Guzmán Zambrano - Juan Pablo Gonzalez Penagos
// Date: 2022-2023
// License: MIT
//
// Description: Builtin definitions
//              (PC port) 
module main

enum __pin_names {    // enumerated type for the pin names
 
    RX=PA11
    TX=PA10


}

fn init() {

}
