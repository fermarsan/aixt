// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Cristian Garzón
// Date: 2023 - 2024
// ## Description
// UART2 functions (WCH-CH573F)

module uart2

fn C.setup(baud_rate u32)
