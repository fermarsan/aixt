module rand

// cstdlib.c
#define     abort(...)              abort(__VA_ARGS__)
#define     srand(...)              srand(__VA_ARGS__)
#define     rand(...)               rand(__VA_ARGS__)
#define     random(...)             Random(__VA_ARGS__)
#define     sys_random_number(...)  SysRandomNumber(__VA_ARGS__)
#define     sys_random_ex(...)      SysRandomEx(__VA_ARGS__)


fn init() {

}