module pin

#define output OUTPUT
#define input INPUT

fn init(){

}