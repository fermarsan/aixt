// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2023-2024
// License: MIT
module uart1

#define uart1__print(MESSAGE)		printf("\033[1;31m");	printf("%s", MESSAGE)	// in red


