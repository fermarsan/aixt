module pin

#define pin.write(PIN, VALUE)	gpio_write(PIN, VALUE)