// Project Name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa - Julian Camilo Guzmán Zambrano - Juan Pablo Gonzalez Penagos
// Date: 2022-2024
// License: MIT
//
// // Description: SLEEP_us functions (Blue-Pill)
//              (PC port) 

module time

#define time__sleep_us(US)    delayMicroseconds(US)