// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2022-2024
// License: MIT
module pin

#define pin__write(PIN_NAME, VALUE) PIN_NAME = VALUE