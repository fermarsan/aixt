module pic16

pub const description = 'API for the PIC16 family devices'
