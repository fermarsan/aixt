module uart

#define uart__setup_1(BAUND_RATE)		Serial1.begin(BAUND_RATE)
