module pwm