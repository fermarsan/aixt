module pin

@[inline]
pub fn write(pin u8, value u8) {
	C.gpio_write(pin, value)
}
