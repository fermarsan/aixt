// Project name: FIRE Hello World
// Author: Fernando M. Santa
// Date: 21/01/2025
// M5Stack FIRE IoT development kit

import lcd
import power

power.setup()	// init the power module
lcd.print("Hello World...")