module uart

fn C.print(msg string)