// Project Name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa - Johann Escobar Guzman - Daniel Andrés Vásquez Gómez
// Date: 2023-2024
// License: MIT
//
// // Description: adc functions (W801)
//              (PC port) 

module pin

#define adc__INPUT   ANALOG_INPUT