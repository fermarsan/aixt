// Author: Fernando M. Santa
// Date: 2025
//
// ## Description
// Builtin definitions (ESP32-DevKitC port)
module main
