module uart

#define uart__println(MESSAGE)   Serial.println(MESSAGE)