// Project Name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa - Johann Escobar Guzmán - Daniel Andrés Vásquez Gómez
// Date: 2023-2024
// License: MIT
//
// // Description: PIN functions (W801)
//              (PC port) 

module pin

#define output		OUTPUT
#define input		INPUT
#define pin__in_pullup	INPUT_PULLUP

fn init() {

}