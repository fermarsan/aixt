module main

fn.init(){

}

