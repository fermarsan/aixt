// Author: Fernando M. Santa
// Date: 2024


// module uart

// // read function reads incoming serial data
// @[as_macro]
// pub fn read_string() string {
// 	return C.SERIAL_READSTRING()
// }
