// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Cristian Garzón
// Date: 2023 - 2024
// ## Description
// UART3 functions (WCH-CH582F)

module uart3

fn C.read() u8
