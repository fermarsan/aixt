module sw_uart

#define sw_uart__setup(BAUDRATE)	sw_uart__baudrate = BAUDRATE