// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: PWM functions (Arduino Mega - ATmega2560 port)
module pwm_fn

@[as_macro] pub const ch0 = 2
@[as_macro] pub const ch1 = 3
@[as_macro] pub const ch2 = 4
@[as_macro] pub const ch3 = 5
@[as_macro] pub const ch4 = 6
@[as_macro] pub const ch5 = 7
@[as_macro] pub const ch6 = 8
@[as_macro] pub const ch7 = 9
@[as_macro] pub const ch8 = 10
@[as_macro] pub const ch9 = 11
@[as_macro] pub const ch10 = 12
@[as_macro] pub const ch11= 13
