// Project Name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: sleep functions (Ai_Thinker_Ai-WB2-32S-Kit)

module time

#define time.sleep(S)    delay(S*1000)