// Project Name: Aixt project, https://gitlab.com/fermarsan/aixt-project.git
// File Name: uart.c.v
// Author: Andrés Felipe Fajardo Duarte and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: UART management functions (PIC18F2550 port)

module uart

#include <xc.h>