// Project name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024-2025
// License: MIT
//
// Description: Builtin definitions
//              (PIC16F676)
module main

#include <xc.h>
#include <stdbool.h>
#include <stdint.h>

#include "builtin.c"


pub fn panic(err string) {

}
