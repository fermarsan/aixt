module time


fn init() {

}