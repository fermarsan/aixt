// Project name: Aixt, https://github.com/fermarsan/aixt.git
//
// _Author:_ Fernando M. Santa
//
// _Date:_ 2025
//
// ## Description
// Aixt's builtin components module
module builtin

// eprint adds a new error message to stderr (Aixt's table error list).
// This function does not generate any code
pub fn eprint(msg string)