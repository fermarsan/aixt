module pwm


fn setup(output u8, freq u16) {
	if output == 1 {
		
	}
}