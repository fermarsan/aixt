module microchip

pub const description = 'API for the Microchip devices'
