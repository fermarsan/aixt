// _File:_ https://github.com/fermarsan/aixt/blob/main/
//
// _Author:_ Fernando M. Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
//
// _Date:_ 2022-2024
//
// // ## Description
// pwm functions (Ai_Thinker_Ai-WB2-32S-Kit)

module pwm

//TODO: add the pin definition
