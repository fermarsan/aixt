// Project Name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa - Daniel Polo - Edwin Barrera
// Date: 2022-2024
// License: MIT
//
// // Description: pin functions (CY8CKIT-049-42XX)

module pin

#define output		OUTPUT
#define input		INPUT
#define in_pullup	INPUT_PULLUP