// Author: Fernando M. Santa - Daniel Polo - Edwin Barrera - Javier Leon - Camilo Lucas
// Date: 2022-2025
//
// ## Description
// pin read functions (CY8CKIT-049-42XX)

module pin

@[as_macro]
pub fn read(name any) u8 {
	return C.PIN_READ(name)
}
