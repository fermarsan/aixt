// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2022-2024
// License: MIT
//
// Description: Builtin definitions (Exp16-PIC24 port)
module main



#include "builtin.c"


// #define led3    A, 0			// Onboard LEDs
// #define led4    A, 1
// #define led5    A, 2
// #define led6    A, 3
// #define led7    A, 4
// #define led8    A, 5
// #define led9    A, 6
// #define led10   A, 7

// #define sw3     D, 6			// Onboard switchs
// #define sw4     D, 13
// #define sw5     A, 7
// #define sw6     D, 7


// fn C.init()