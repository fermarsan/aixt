module uart2

fn C.write(data u8)