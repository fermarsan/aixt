module pic12

pub const description = 'API for the PIC12 family devices'
