module pic16f8x

pub const description = 'API for the PIC16F8x family devices'
