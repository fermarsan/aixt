module main

#include "CH58x_common.h"

fn init() {
	// SetSysClock(CLK_SOURCE_PLL_60MHz)
}
