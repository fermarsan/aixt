// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: PWM functions W801
module pwm

pub const ch0_0 = u8(C.PA2)
pub const ch0_1 = u8(C.PA10)
pub const ch0_2 = u8(C.PB0)
pub const ch0_3 = u8(C.PB12)
pub const ch0_4 = u8(C.PB19)

pub const ch1_0 = u8(C.PA3)
pub const ch1_1 = u8(C.PA11)
pub const ch1_2 = u8(C.PB1)
pub const ch1_3 = u8(C.PB13)
pub const ch1_4 = u8(C.PB20)

pub const ch2_0 = u8(C.PA0)
pub const ch2_1 = u8(C.PA12)
pub const ch2_2 = u8(C.PB2)
pub const ch2_3 = u8(C.PB14)
pub const ch2_4 = u8(C.PB24)

pub const ch3_0 = u8(C.PA1)
pub const ch3_1 = u8(C.PA13)
pub const ch3_2 = u8(C.PB3)
pub const ch3_3 = u8(C.PB15)
pub const ch3_4 = u8(C.PB25)

pub const ch4_0 = u8(C.PA4)
pub const ch4_1 = u8(C.PA7)
pub const ch4_2 = u8(C.PA14)
pub const ch4_3 = u8(C.PB16)
pub const ch4_4 = u8(C.PB26)