module Microchip

pub const description = 'Workspace for the Microchip devices'
