module string

// cstring.h
#define     string__to_num(...)              StrToNum(__VA_ARGS__)
#define     string__str_len(...)             StrLen(__VA_ARGS__)
#define     string__index(...)               StrIndex(__VA_ARGS__)
#define     string__num_to(...)              NumToStr(__VA_ARGS__)
#define     string__str_cat(...)             StrCat(__VA_ARGS__)
#define     string__sub(...)                 SubStr(__VA_ARGS__)
#define     string__flatten(...)             Flatten(__VA_ARGS__)
#define     string__replace(...)             StrReplace(__VA_ARGS__)
#define     string__format_num(...)          FormatNum(__VA_ARGS__)
#define     string__format_val(...)          FormatVal(__VA_ARGS__)
#define     string__flatten_var(...)         FlattenVar(__VA_ARGS__)
#define     string__unflatten_var(...)       UnflattenVar(__VA_ARGS__)
#define     string__pos(...)                 Pos(__VA_ARGS__)
#define     string__byte_array_to(...)       ByteArrayToStr(__VA_ARGS__)
#define     string__byte_array_to_ex(...)    ByteArrayToStrEx(__VA_ARGS__)
#define     string__to_byte_array(...)       StrToByteArray(__VA_ARGS__)
#define     string__copy(...)                Copy(__VA_ARGS__)
#define     string__mid(...)                 MidStr(__VA_ARGS__)
#define     string__right(...)               RightStr(__VA_ARGS__)
#define     string__left(...)                LeftStr(__VA_ARGS__)
#define     string__len(...)                 strlen(__VA_ARGS__)
#define     string__cat(...)                 strcat(__VA_ARGS__)
#define     string__n_cat(...)               strncat(__VA_ARGS__)
#define     string__cpy(...)                 strcpy(__VA_ARGS__)
#define     string__n_cpy(...)               strncpy(__VA_ARGS__)
#define     string__cmp(...)                 strcmp(__VA_ARGS__)
#define     string__n_cmp(...)               strncmp(__VA_ARGS__)
#define     string__memcpy(...)              memcpy(__VA_ARGS__)
#define     string__memmove(...)             memmove(__VA_ARGS__)
#define     string__memcmp(...)              memcmp(__VA_ARGS__)
#define     string__address_of(...)          addressOf(__VA_ARGS__)
#define     string__reladdress_of(...)       reladdressOf(__VA_ARGS__)
#define     string__address_of_ex(...)       addressOfEx(__VA_ARGS__)

// Functions for use with NXC array types.
#define		string__upper_case(...) 	UpperCase(__VA_ARGS__) 
#define		string__lower_case(...) 	LowerCase(__VA_ARGS__) 
#define		string__upper_case_ex(...) 	UpperCaseEx(__VA_ARGS__) 
#define		string__lower_case_ex(...) 	LowerCaseEx(__VA_ARGS__) 
