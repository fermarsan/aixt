// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2023-2024
// License: MIT
//
// Description: This is a module to emulate ADC inputs in console.
module adc

// Channel_names is the enumerated type for the ADC channel names
enum Channel_names {
    ch_0 = 0
    ch_1   
}

__global (
    value__ = 0
)

fn init() {
    
}