// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: 
// Date: 
// License: MIT
//
// Description: 
module port

#define TRISa	TRISA	// port setup name equivalents
#define TRISb	TRISB
...

#define PORTa	PORTA	// port in name equivalents
#define PORTb	PORTB
...

#define LATa	LATA	// port out name equivalents (PIC18, PIC24, dsPIC33)
#define LATb	LATB	
...
