// Project Name: Aixt, https://github.com/fermarsan/aixt.git

// Author: Jan Carlo Peñuela Jurado and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: ADC
//              (PIC18F452)
module adc
#include <xc.h>

fn init() {
    
}