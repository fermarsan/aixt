// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Authors:
//		- Jahn Delgado
//		- Fernando M. Santa
// Date: 22/05/2025
// License: MIT
//
// Description: Builtin definitions (ESP32-CYD 2.8 inch)
//
module main
