// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: high.c.v
// Author: Fernando Martínez Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: HIGH functions (Ai_Thinker_Ai-WB2-32S-Kit)

module pin

#define pin__high(PIN_NAME)   digitalWrite(PIN_NAME, HIGH)