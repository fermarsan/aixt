module main



