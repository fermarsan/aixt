module pwm

#define pwm__write(PIN, VAL)	analogWrite(PIN, VAL)
