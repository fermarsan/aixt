module nano

pub const description = 'Arduino Nano target API'
