// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: pin.c.v
// Author: Fernando M. Santa - Johann Escobar Guzmán - Daniel Andrés Vásquez Gómez
// Date: 2023-2024
// License: MIT
//
// // Description: PIN functions (W801)
//              (PC port) 

module pin

#define pin__output		OUTPUT
#define pin__input		INPUT
#define pin__in_pullup	INPUT_PULLUP

fn init() {

}