// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// File Name: pwm.c.v
// Author: Andrés Felipe Fajardo Duarte and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: PWM management functions (PIC18F2550 port)

module pwm 

#include <xc.h>

fn init() {
    
}