// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git
// File Name: read.c.v
// Author: Fernando Martinez Santa - Arley Junco - Luis Quevedo 
// Date: 2024
// License : MIT

module pin 

#define pin_read(PIN_NAME)   digitalRead(PIN_NAME)