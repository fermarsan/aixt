module avr

pub const description = 'Arduino AVR based devices API'
