module pic16f6xx_20p

pub const description = 'API for the PIC16f6xx_20p family devices'
