// Project Name : Aixt: http://github.com/fermansan/aixt.git
//
// _Author:_ Farith Ochoa León, Delipe Cardozo and Fernando M. Santa 
// License : MIT
//
// _Date:_ 2024-2025

module pwm 


@[as_macro] pub const ch0 = 0 
@[as_macro] pub const ch1 = 1
@[as_macro] pub const ch2 = 2
@[as_macro] pub const ch3 = 3
@[as_macro] pub const ch4 = 4
@[as_macro] pub const ch5 = 5
@[as_macro] pub const ch6 = 6
@[as_macro] pub const ch7 = 7
@[as_macro] pub const ch8 = 8
@[as_macro] pub const ch9 = 9
@[as_macro] pub const ch10 = 10

@[as_macro] pub const ch18 = 18
@[as_macro] pub const ch19 = 19
@[as_macro] pub const ch20 = 20
@[as_macro] pub const ch21 = 21