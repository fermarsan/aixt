// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git
// File Name: uart.c.v
// Author: Farith Ochoa Leon, Felipe Cardozo and Fernando Martinez Santa
// Date: 2024
// License : MIT

module uart 

fn init() {
	
}