module uart

fn init(){

}