// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: dutymax.c.v
// Author: Fernando Martínez Santa - Johann Escobar Guzmán - Daniel Andrés Vásquez Gómez
// Date: 2023-2024
// License: MIT
//
// // Description: DUTY_MAX functions (W801)
//              (PC port) 

module pin

#define DUTY__MAX  DUTY_MAX