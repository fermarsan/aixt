// Project Name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa - Johann Escobar Guzman - Daniel Andrés Vásquez Gómez
// Date: 2024
// License: MIT
//
// Description: ADC management functions (W801)
module adc

fn C.setup(pins u16, fad u8, nbits u8)