module nxt

pub const description = 'API for the Mindstorms NXT target'
