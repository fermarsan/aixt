// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2022-2024
// License: MIT
module pin

#define pin__setup(PIN_NAME, PIN_MODE)   PIN_NAME = PIN_MODE
