module pin

#define pin__setup(PIN_NUMBER, PIN_MODE)	printf("TRIS ## PIN_NUMBER ## bits.TRIS ## PIN_NUMBER = PIN_MODE")