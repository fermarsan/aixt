module adc

  adc__setup(PIN_NAME, SETUP_VALUE)
