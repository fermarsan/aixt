// Project Name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: setup functions (Ai_Thinker_Ai-WB2-32S-Kit)

module pin

#define pin.setup(PIN_NAME, MODE)    pinMode(PIN_NAME, MODE)