// Author: Fernando M. Santa
// Date: 2024
//
// ## Description
// ADC functions
module adc2

// adc channels
pub const ch0 = 4
pub const ch1 = 0
pub const ch2 = 2
pub const ch3 = 15
pub const ch4 = 13
pub const ch5 = 12
pub const ch6 = 14
pub const ch7 = 27
// pub const ch8 = xx
pub const ch9 = 26