// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: adcinput.v
// Author: Fernando Martínez Santa - Johann Escobar Guzman - Daniel Andrés Vásquez Gómez
// Date: 2023-2024
// License: MIT
//
// // Description: adc functions (W801)
//              (PC port) 

module pin

#define adc__INPUT   ANALOG_INPUT