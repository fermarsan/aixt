// Project name: Aixt, https://github.com/fermarsan/aixt.git
//
// _Author:_ Fernando M. Santa
//
// _Date:_ 2025
// License: MIT
module pin

#include "toggle.c"

fn C.DIGITAL_TOGGLE(id u8)

// toggle function toggles the value to a specific pin
// @[as_macro]
@[inline]
pub fn (mut p Pin) toggle() {   
    C.DIGITAL_TOGGLE(p.id)
}