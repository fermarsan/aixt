module uart2

fn C.setup(baud_rate u32)