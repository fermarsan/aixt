// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
//
// ## Description
// PWM functions (Arduino Uno - ATmega328P port)
module pwm

@[as_macro] pub const ch0 = 3
@[as_macro] pub const ch1 = 5
@[as_macro] pub const ch2 = 6
@[as_macro] pub const ch3 = 9
@[as_macro] pub const ch4 = 10
@[as_macro] pub const ch5 = 11
