// File: https://github.com/fermarsan/aixt/blob/main/
// Author: Fernando M. Santa - Daniel Polo - Edwin Barrera - Javier Leon - Camilo Lucas
// Date: 2022-2025
//
// // ## Description
// low functions (CY8CKIT-145-40XX)



module pin

@[as_macro]
pub fn low(name any) {
	C.PIN_LOW(name)
}
