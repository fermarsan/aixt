module pin

#define pin__out OUTPUT
#define pin__in INPUT
fn.init(){

}