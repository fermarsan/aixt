module pwm
fn_init(){

}