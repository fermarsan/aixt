// Project Name : Aixt: http://github.com/fermansan/aixt.git
//
// _Author:_ Fernando M. Santa 
// License : MIT
//
// _Date:_ 2025

module pwm 


pub const ch0 = 0 
pub const ch1 = 1
pub const ch2 = 2
pub const ch3 = 3
pub const ch4 = 4
pub const ch5 = 5
pub const ch6 = 6
pub const ch7 = 7
pub const ch8 = 8
pub const ch9 = 9
pub const ch10 = 10
pub const ch11 = 11
pub const ch12 = 12
pub const ch13 = 13

pub const ch18 = 18
pub const ch19 = 19