// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Pin management functions Arduino devices
module pin

// pin names
pub const gp0   = 0    
pub const gp1   = 1
pub const gp2   = 2
pub const gp3   = 3
pub const gp4   = 4
pub const gp5   = 5
pub const gp6   = 6
pub const gp7   = 7
pub const gp8   = 8
pub const gp9   = 9
pub const gp10  = 10
pub const gp11  = 11
pub const gp12  = 12
pub const gp13  = 13
pub const gp14  = 14
pub const gp15  = 15
pub const gp16  = 16
pub const gp17  = 17
pub const gp18  = 18
pub const gp19  = 19
pub const gp20  = 20
pub const gp21  = 21
pub const gp22  = 22
pub const _gp23 = 23
pub const _gp24 = 24
pub const gp25  = 25
pub const gp26  = 26
pub const gp27  = 27
pub const gp28  = 28
