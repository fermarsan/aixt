// Project Name : Aixt: http://github.com/fermansan/aixt.git
//
// _Author:_ Farith Ochoa León, Delipe Cardozo and Fernando M. Santa 
// License : MIT
//
// _Date:_ 2024-2025
//
// ## Description
// ADC functions
module adc2

// ADC pin names
pub const ch0 = 5