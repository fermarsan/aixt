module main

#include "CH82x_common.h"
#define true 1

//fn init() {
	//SetSysClock(CLK_SOURCE_PLL_60MHz)
//}
