// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: builtin.c
// Author: Fernando Martínez Santa - Julian Camilo Guzmán Zambrano - Juan Pablo Gonzalez Penagos
// Date: 2022-2023
// License: MIT
//
// Description: Builtin definitions
//              (PC port) 
module main

enum __pin_names {    // enumerated type for the pin names
 
    rX=PA11
    tX=PA10
    p1=PA0
    p2=PA1
    p3=PA2
    p4=PA3
    p5=PA4
    p6=PA5
    p7=PA6
    p8=PA7
    p9=PB0
    p10=PB1
    p11=PB10
    p12=PB11
    p13=PB12
    p14=PB13
    p15=PB14
    p16=PB15
    p17=PA8
    p18=PB3
    p19=PB4
    p20=PB5
    p21=PB6
    p22=PB7
    p23=PB8
    p24=PB9
    p25=PC13
    recibe_dato
    dato
    envia_dato

}

fn init() {

}
