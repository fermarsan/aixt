// Project Name: Aixt project, https://gitlab.com/fermarsan/aixt-project.git
// File Name: time.c.v
// Author: Jan Carlo Peñuela Jurado and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: TIME function
//              (PIC18F452)


module time

#include <xc.h>