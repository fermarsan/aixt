module time

#define time.sleep_ms(MS)    delay(MS)