// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Cristian Garzón
// Date: 2023 - 2024
// Description: TIME functions (WCH-CH582F)

module time

#define time.sleep_ms(TIME)    DelayMs(TIME)

