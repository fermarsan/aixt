// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fabián A. Rojas Acosta, Alberto Pinzón Valero and Fernando M. Santa
// Date: 2024
// License: MIT
module time

//Pauses the program for the amount of time (in seconds) specified as parameter
#define time.sleep(TS)  delay(TS*1000)