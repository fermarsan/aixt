// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git

// Author: Fernando M. Santa - Arley Junco - Luis Quevedo 
// Date: 2024
// License : MIT

module uart 

#define TX_PIN PD6
#include "ATtinySerialOut.hpp"

fn init() {
	
}