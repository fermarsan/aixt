// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Cristian Garzón
// Date: 2023 - 2024
// Description: PWM functions (WCH-CH573F)

module pwm

/* CHANNEL 4  PIN A12
   CHANNEL 5  PIN A13
   CHANNEL 7  PIN B4 
   CHANNEL 9  PIN B7 
   CHANNEL 10 PIN B14
   CHANNEL 11 PIN 23 */ 

   