module pin

#define pin.write(PIN_NAME, VALUE)		digitalWrite(PIN_NAME, VALUE)
