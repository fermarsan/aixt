module math

const (
	pi = 3.141592
	e = 2.71828
)