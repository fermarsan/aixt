// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 29/01/2025
// License: MIT
//
// Description: Example of a Library module.
//
module ex_array

fn C.ArrayMin(src []any, idx u16, len u16) any