module uart
#define uart__Write(VALUE)    Serial.write(VALUE)