module pin

#define pin.read(PIN_NAME)		digitalRead(PIN_NAME)
