module time


