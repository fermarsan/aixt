// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: pin.c.v
// Author: Fernando Martínez Santa - Julian Camilo Guzmán Zambrano - Juan Pablo Gonzalez Penagos
// Date: 2022-2024
// License: MIT
//
// // Description: PIN functions (Blue Pill_STM32F103C)
//              (PC port) 

module pin

#define pin__output		OUTPUT
#define pin__input			INPUT
#define pin__in_pullup	INPUT_PULLUP

fn init() {

}