module uart2

