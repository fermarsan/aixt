module pin

#define output		OUTPUT
#define input		INPUT
#define pin__in_pullup	INPUT_PULLUP

fn init() {

}