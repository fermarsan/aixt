module uart2

fn C.print(msg string)