// Author: Cesar Alejandro Roa Acosta and Fernando M. Santa
// Date: 2024-2025
//
// ## Description
// Builtin definitions
//              (PIC16F87x)
module main

#include <xc.h>
#include <stdbool.h>
#include <stdint.h>

#include "main.c"
