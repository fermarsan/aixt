// Project Name : Aixt: http://github.com/fermansan/aixt.git
// Author: Farith Ochoa León, Delipe Cardozo and Fernando M. Santa 
// License : MIT

module pin 

#define output 		OUTPUT 
#define input 			INPUT
#define input_pullup 	INPUT_PULLUP

fn init () { 
	
}