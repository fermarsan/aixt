module pin

#define pin__setup(PIN,  MODE)   gpio_set_mode(PIN, MODE)