// _File:_ https://github.com/fermarsan/aixt/blob/main/
// Authors:
//	 - Julian Camilo Guzmán Zambrano
//	 - Juan Pablo Gonzalez Penagos
//	 - Fernando M. Santa
//
// _Date:_ 2022-2025
//
// ## Description
// Builtin definitions (Blue-Pill port)
module main
