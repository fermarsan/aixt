// Project Name: Aixt project, https://gitlab.com/fermarsan/aixt-project.git
// File Name: builtin.c.v
// Author: Farith Ochoa León and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: Builtin definitions (ESP32-C3FH4)
//              

module main

fn init() { 

}
