// Author: Fernando M. Santa - Daniel Polo - Edwin Barrera - Javier Leon - Camilo Lucas
// Date: 2022-2025
//
// ## Description
// pin functions (CY8CKIT-145-40XX)

module pin

#include "pin.c"


fn C.PIN_WRITE(name any, value any)
fn C.PIN_HIGH(name any)
fn C.PIN_LOW(name any)
fn C.PIN_READ(name any) u8
