// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024-2025
// License: MIT
//
// Description: ADC functions
module adc

fn C.analogReadResolution(res any)

// adc channels
pub const ch0 = u8(C.A0)
pub const ch1 = u8(C.A1)
pub const ch2 = u8(C.A2)
pub const ch3 = u8(C.A3)
pub const ch4 = u8(C.A4)
pub const ch5 = u8(C.A5)
pub const ch6 = u8(C.A6)
pub const ch7 = u8(C.A7)
pub const ch8 = u8(C.A8)
pub const ch9 = u8(C.A9)
pub const ch10 = u8(C.A10)
