// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2023-2024
// License: MIT
//
// Description: This is a module to emulate ADC inputs in console.
module adc

enum ADC_names {
    an0 = 0
    ch1      
}