// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Jan Carlo Peñuela y Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Pin port management functions (PIC18F2550 port)

module port

#include <xc.h>

const output = C.0   // port mode (direction)
const input = C.1


