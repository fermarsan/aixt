// Project Name: Aixt project, https://gitlab.com/fermarsan/aixt-project.git
// File Name: port.c.v
// Author: Luis Alfredo Pinto Medina and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: Pin-port functions (PIC16F84A port)

module port

#define TRISa	TRISA	// port setup name equivalents
#define TRISb	TRISB
#define TRISc	TRISC
#define TRISd	TRISD
#define TRISe	TRISE
#define TRISf	TRISF
#define TRISg	TRISG

#define PORTa	PORTA	// port in name equivalents
#define PORTb	PORTB
#define PORTc	PORTC
#define PORTd	PORTD
#define PORTe	PORTE
#define PORTf	PORTF
#define PORTg	PORTG

