// Author: Fernando M. Santa
// Date: 29/01/2025
//
// ## Description
// Example of a Library module.
//
module ex_array

fn C.min(a any, b any) any