module pwm


fn C.setup(output u8, freq u16) 