// Project Name: Aixt project, https://gitlab.com/fermarsan/aixt-project.git
// File Name: time.c.v
// Author: Luis Alfredo Pinto Medina and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: seconds delay function
//              (PIC16F886 port)

module time

fn init() {

}