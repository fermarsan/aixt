// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2023-2024
// License: MIT
//
// Description: This is a module to emulate ADC inputs in console.
module adc

pub const (
    ch0 = 0   // adc channel
    ch1 = 1   // constants
)