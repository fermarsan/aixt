// module importing

import time { sleep }
import machine

a := 0

for {
	sleep(1000)
	a++
}