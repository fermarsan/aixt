// Project name: Aixt, https://github.com/fermarsan/aixt.git
//
// _Author:_ Cristian Garzón
//
// _Date:_ 2023 - 2024
// ## Description
// UART functions (WCH-CH573F)

module uart

fn C.setup(baud_rate u32)
