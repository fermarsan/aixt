module math

// Miscellaneous NBC/NXC constants
#define 	math__pi					  PI
#define 	math__rad_to_deg			  RADIANS_PER_DEGREE
#define 	math__deg_to_rad			  DEGREES_PER_RADIAN

// cmath.h
#define     math__sqrt(...)               sqrt(__VA_ARGS__)
#define     math__cos(...)                cos(__VA_ARGS__)
#define     math__sin(...)                sin(__VA_ARGS__)
#define     math__tan(...)                tan(__VA_ARGS__)
#define     math__acos(...)               acos(__VA_ARGS__)
#define     math__asin(...)               asin(__VA_ARGS__)
#define     math__atan(...)               atan(__VA_ARGS__)
#define     math__atan2(...)              atan2(__VA_ARGS__)
#define     math__cosh(...)               cosh(__VA_ARGS__)
#define     math__sinh(...)               sinh(__VA_ARGS__)
#define     math__tanh(...)               tanh(__VA_ARGS__)
#define     math__exp(...)                exp(__VA_ARGS__)
#define     math__log(...)                log(__VA_ARGS__)
#define     math__log10(...)              log10(__VA_ARGS__)
#define     math__trunc(...)              trunc(__VA_ARGS__)
#define     math__frac(...)               frac(__VA_ARGS__)
#define     math__pow(...)                pow(__VA_ARGS__)
#define     math__ceil(...)               ceil(__VA_ARGS__)
#define     math__floor(...)              floor(__VA_ARGS__)
#define     math__muldiv32(...)           muldiv32(__VA_ARGS__)
#define     math__cosd(...)               cosd(__VA_ARGS__)
#define     math__sind(...)               sind(__VA_ARGS__)
#define     math__tand(...)               tand(__VA_ARGS__)
#define     math__acosd(...)              acosd(__VA_ARGS__)
#define     math__asind(...)              asind(__VA_ARGS__)
#define     math__atand(...)              atand(__VA_ARGS__)
#define     math__atan2d(...)             atan2d(__VA_ARGS__)
#define     math__coshd(...)              coshd(__VA_ARGS__)
#define     math__sinhd(...)              sinhd(__VA_ARGS__)
#define     math__tanhd(...)              tanhd(__VA_ARGS__)
#define     math__bcd2dec(...)            bcd2dec(__VA_ARGS__)
#define     math__is_nan(...)             isNAN(__VA_ARGS__)
#define     math__sign(...)               sign(__VA_ARGS__)
#define     math__vector_cross(...)       VectorCross(__VA_ARGS__)
#define     math__vector_dot(...)         VectorDot(__VA_ARGS__)
#define     math__vector_normalize(...)   VectorNormalize(__VA_ARGS__)

// cstdlib.c
#define     math__abs(...)                abs(__VA_ARGS__)
#define     math__labs(...)               labs(__VA_ARGS__)
#define     math__div(...)                div(__VA_ARGS__)
#define     math__ldiv(...)               ldiv(__VA_ARGS__)


fn init() {
	
}