// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: read.c.v
// Author: Fernando Martínez Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: READ functions (Ai_Thinker_Ai-WB2-32S-Kit)
//              (PC port) 

module pin

#define pin__read(PIN_NAME)   digitalRead(PIN_NAME)