module uart
fn.init(){

}