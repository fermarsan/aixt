// Author: Fernando M. Santa
// Date: 2022-2024
//
// ## Description
// Builtin definitions (Exp16-PIC24 port)
module main

#include <xc.h>
#include <stdint.h>
#include <stdbool.h>

#include "main.c"




// fn C.init()
