// Project Name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Pin-port functions (PIC16F8x port)
module port

enum Port__names as u8 {
	port__a = 0
	port__b
	port__c
	port__d
	port__e 
}
