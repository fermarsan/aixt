// File: https://github.com/fermarsan/aixt/blob/main/
// Author: Fernando M. Santa
// Date: 2022-2025
//
// ## Description
// Builtin definitions (XIAO-SAMD21 port)
module main
