// File: https://github.com/fermarsan/aixt/blob/main/
// Authors:
//	- Luis Alfredo Pinto Medina
//	- Fernando M. Santa
// Date: 2024
//
// ## Description
// Builtin definitions (PIC16F8x port)

module main

#include <xc.h>
#include <stdint.h>
#include <stdbool.h>

#include "builtin.c"
