module ui

// 