module uart

#define	uart__any()	U1STAbits.URXDA