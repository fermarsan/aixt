// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: builtin.c.v
// Author: Fernando Martínez Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: Builtin definitions

module main

enum __pin_names {    // enumerated type for the pin names
    io11=11
    io14=14
    io17=17
    io3=3
    io4=4
    io5=5
    io7=7
    io16=16
    io12=12
}

fn init() {

}
