// Project Name: Aixt project, https://gitlab.com/fermarsan/aixt-project.git
// File Name: port.c.v
// Author: Cesar Alejandro Roa Acosta and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: Port management functions
//              (PIC16F676 port)

module port

fn init() {
    
}