module adc

fn init() {
	
}