// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Builtin definitions (Arduino Mega - ATmega2560 port)
module main


@[as_macro]	const led_0 = 13
