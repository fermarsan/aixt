module pwm

#define pwm__write(PIN_NAME, MODE)   analogWrite(PIN_NAME, MODE)
