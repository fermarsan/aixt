// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Time module (Arduino devices)
module time


fn C.delay(tms int)
fn C.delayMicroseconds(tus int)