module uart

fn init() {

}