// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Pin management functions Arduino devices
module pin

// pin names
pub const gpio0 = 0      
pub const gpio1 = 1  
pub const gpio2 = 2  
pub const gpio3 = 3  
pub const gpio4 = 4  
pub const gpio5 = 5  
pub const gpio6 = 6  
pub const gpio7 = 7  
pub const gpio8 = 8  
pub const gpio9 = 9  
pub const gpio10 = 10   
pub const gpio11 = 11   
pub const gpio12 = 12   
pub const gpio13 = 13   
pub const gpio14 = 14   
pub const gpio15 = 15   
pub const gpio16 = 16   
pub const gpio17 = 17   
pub const gpio18 = 18   
pub const gpio19 = 19   
pub const gpio20 = 20   
pub const gpio21 = 21   
pub const gpio22 = 22   
pub const gpio23 = 23   
pub const gpio24 = 24   
pub const gpio25 = 25   
pub const gpio26 = 26   
pub const gpio27 = 27   
pub const gpio28 = 28   
pub const gpio29 = 29 
pub const gpio30 = 30 
pub const gpio31 = 31 
pub const gpio32 = 32 
pub const gpio33 = 33 
pub const gpio34 = 34 
pub const gpio35 = 35 
pub const gpio36 = 36 
pub const gpio39 = 39

// pin modes
pub const input		= u8(C.INPUT)
pub const output	= u8(C.OUTPUT)
pub const in_pullup = u8(C.INPUT_PULLUP)

