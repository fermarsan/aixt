// Project Name: Aixt project, https://gitlab.com/fermarsan/aixt-project.git
// File Name: Digital.c.v
// Author: Cesar Alejandro Roa Acosta and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: Digital management functions
//              (PIC16F676 port)

module pin 

#define pin__digital()  ANSEL = 0

