module uart

#define uart__println_1(MESSAGE)   Serial1.println(MESSAGE)