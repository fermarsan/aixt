// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: 
//	- Fabián A. Rojas Acosta
//	- Alberto Pinzón Valero
//	- Fernando M. Santa
// Date: 2024-2025
// License: MIT
//
// Description: Builtin definitions (Arduino Nano - ATmega328P port)
module main

#include "builtin.c"
