// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2023-2024
// License: MIT
module uart2

#define uart2__print(MESSAGE)		printf("\033[1;34m");	printf("%s", MESSAGE)	// in blue

