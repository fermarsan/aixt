module pin

#define pin.setup(PIN,  MODE)   gpio_set_mode(PIN, MODE)