module pwm

#define pwm.write(PIN, VAL)	analogWrite(PIN, VAL)