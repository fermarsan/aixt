// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// File Name: pwm.c.v
// Author: Jan Carlo Peñuela Jurado and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: PWM
//              (PIC18F452)
module pwm
#include <xc.h>

fn init() {
    
}