// Project Name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa - Johann Escobar Guzmán - Daniel Andrés Vásquez Gómez
// Date: 2023-2024
// License: MIT
//
// // Description: SLEEP_ms functions (W801)
//              (PC port) 

module uart

#define uart.print_0(MESSAGE)	Serial.print(MESSAGE)

#define uart.print_1(MESSAGE)	Serial1.print(MESSAGE)

#define uart.print_x(UART_NUMBER, MESSAGE)		uart.print_ ## UART_NUMBER (MESSAGE) 			

// macro with 1 or 2 arguments
#define SEL_uart.print(_1, _2, MACRO_NAME, ...) MACRO_NAME
#define uart.print(...) SEL_uart.print(__VA_ARGS__, uart.print_x, uart.print_0)(__VA_ARGS__)