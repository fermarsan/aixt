// Project Name : Aixt: http://github.com/fermansan/aixt.git
// Authors:
//	- Farith Ochoa Leon
//	- Felipe Cardozo
//	- Fernando M. Santa
// Date: 2024-2025
// License : MIT
//
//Description: Builtin definitions (ESP32-C3FH4)      

module main

// builtin LED
const led_0 = u8(12)
const led_1 = u8(13)

