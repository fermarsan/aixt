// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: ready_1.c.v
// Author: Fernando Martínez Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: READY_1 functions (Ai_Thinker_Ai-WB2-32S-Kit)
//              (PC port) 

module uart

#define uart__ready_1   Serial1.available