// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fabián A. Rojas Acosta, Alberto Pinzón Valero and Fernando Martínez Santa
// Date: 2024
// License: MIT
module time

//Pauses the program for the amount of time (in milliseconds) specified as parameter
#define time__sleep_ms(TMS)  delay(TMS)