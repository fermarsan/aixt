// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git
// File Name: pwm.c.v
// Author: Fernando Martinez Santa - Arley Junco - Luis Quevedo 
// Date: 2024
// License : MIT

module pwm

fn init() {
	
}