module main

fn init() {
	
}