// Project Name : Aixt: http://github.com/fermansan/aixt.git
// Author: Farith Ochoa León, Delipe Cardozo and Fernando M. Santa 
// License : MIT
// Date: 2024-2025
//
// Description: ADC functions
module adc

// ADC pin names
@[as_macro] pub const ch0 = 0
@[as_macro] pub const ch1 = 1
@[as_macro] pub const ch2 = 2
@[as_macro] pub const ch3 = 3
@[as_macro] pub const ch4 = 4
@[as_macro] pub const ch5 = 5