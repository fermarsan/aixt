// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git
// File Name: low.c.v
// Author: Fernando M. Santa - Arley Junco - Luis Quevedo 
// Date: 2024
// License : MIT

module pin

#define pin__low(PIN_NAME)        digitalWrite(PIN_NAME, LOW)