module adc
