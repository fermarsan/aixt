// Project name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Cesar Alejandro Roa Acosta and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Port management functions
//              (PIC16F676 port)
module port

#define TRISa		TRISA	// port setup name equivalents
#define TRISc		TRISC

#define PORTa		PORTA	// port in name equivalents
#define PORTc		PORTC