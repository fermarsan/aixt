module time
fn.init(){

}
