module uart

fn C.setup(baud_rate u32)