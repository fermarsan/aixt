// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Builtin definitions (Arduino Mega - ATmega2560 port)
module main

#include "builtin.c"

// builtin LED
@[as_macro]	const led0 = 13