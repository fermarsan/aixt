module main


