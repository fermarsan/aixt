// Author: Fernando M. Santa
// Date: 2024-2025
//
// ## Description
// Builtin definitions
//              (PIC16F676)
module main

#include <xc.h>
#include <stdbool.h>
#include <stdint.h>

#include "main.c"
