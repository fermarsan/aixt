module pwm

#define pwm_write(PIN_NAME, MODE)   analogWrite(PIN_NAME, MODE)