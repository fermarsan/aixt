module time

fn init() {

}
