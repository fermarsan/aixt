// Project Name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa - Johann Escobar Guzmán - Daniel Andrés Vásquez Gómez
// Date: 2023-2024
// License: MIT
//
// // Description: PIN functions (W801)
//              (PC port) 

module pin
#define pwm.pin[PIN_NAME]  pwm_pin[PIN_NAME]