// Project Name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa - Daniel Polo - Edwin Barrera
// Date: 2022-2024
// License: MIT
//
// // Description: pin functions (CY8CKIT-145-40XX)

module pin

#include "pin.c"


fn C.PIN_WRITE(name any, value any) 