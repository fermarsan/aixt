module pin

#define pin__output OUTPUT
#define pin__input INPUT

