module time

#define time__sleep_ms(TIME)	mtimer_delay_ms(TIME)