module time

#define time__sleep_ms(TIME)  delay(TIME)
fn_init(){

}