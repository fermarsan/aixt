module uart

