// Project Name: Aixt project, https://gitlab.com/fermarsan/aixt-project.git
// File Name: builtin.c.v
// Author: Farith Ochoa León, Felipe Cardozo Hernandez and Fernando Martínez Santa
// Date: 2024
// License: MIT

module time

#define time__sleep_ms(TIME)      delay(TIME)