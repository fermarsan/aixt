// Project Name : Aixt: http://github.com/fermansan/aixt.git
// Author: Farith Ochoa León, Delipe Cardozo and Fernando M. Santa 
// License : MIT

module adc 

@[inline]
pub fn read(PIN_NAME) {
C.analogRead(PIN_NAME)
}
