module uart

#define uart__setup_1(BAUD_RATE)   Serial1.begin(BAUD_RATE)