// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git
// File Name: time.c.v
// Author: Fernando Martinez Santa - Arley Junco - Luis Quevedo 
// Date: 2024
// License : MIT

module time

fn init() {
	
}