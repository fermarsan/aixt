module adc

#define adc.read(PIN_NAME)   analogRead(PIN_NAME)