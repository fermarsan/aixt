module uart2

fn C.read() u8