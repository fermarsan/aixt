// Project Name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: Pin-port functions (ATmega328p)
module port

enum Port__names as u8 {
	port__b = 0
	port__c
	port__d
}
