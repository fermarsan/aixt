// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024-2025
// License: MIT
//
// Description: ADC functions
module adc

// adc channels
pub const ch0 = u8(C.A0)
pub const ch1 = u8(C.A1)
pub const ch2 = u8(C.A2)