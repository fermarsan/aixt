
module pin

#define pin.setup(PIN_NAME, MODE)    pinMode(PIN_NAME, MODE)