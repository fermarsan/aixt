// _File:_ https://github.com/fermarsan/aixt/blob/main/
//
// _Author:_ Fernando M. Santa
//
// _Date:_ 2022-2025
//
// ## Description
// Builtin definitions (Nucleo-L031K6 port)
module main

// builtin LED
const led0 = 13
