// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Authors:
//		- Jahn Delgado
//		- Fernando M. Santa
//
// _Date:_ 22/05/2025
//
// ## Description
// Builtin definitions (ESP32-CYD 2.8 inch)
//
module main
