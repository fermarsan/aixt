// Project Name : Aixt: http://github.com/fermansan/aixt.git
// Authors:
//  - Arley Junco
//  - Luis Quevedo
//  - Fernando M. Santa
// Date: 2024
// License : MIT


module pin

#  define output 			OUTPUT
#  define input  			INPUT  
#  define input_pullup  	INPUT_PULLUP

