// _File:_ https://github.com/fermarsan/aixt/blob/main/
//
// _Author:_ Fernando M. Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
//
// _Date:_ 2022-2024
//
// // ## Description
// Builtin definitions

module main
