module uart

#define uart__read()		Serial.read()
