// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git

// Author: Fernando M. Santa - Arley Junco - Luis Quevedo 
// Date: 2024
// License : MIT


module pin

# define pin__output 			OUTPUT
# define pin__input  			INPUT  
# define pin__input_pullup  	INPUT_PULLUP

fn init() {

}