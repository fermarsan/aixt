module pin

#define pin__low(PIN_NAME)		digitalWrite(PIN_NAME, LOW)
fn.init(){

}