// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git

// Author: Farith Ochoa León, Delipe Cardozo and Fernando M. Santa 
// License : MIT

module pin 

#define output 		OUTPUT 
#define input 			INPUT
#define input_pullup 	INPUT_PULLUP

fn init () { 
	
}