// Author: Fernando M. Santa
// Date: 2022-2025
//
// ## Description
// Builtin definitions (Nucleo-L031K6 port)
module main

// builtin LED
const led0 = 13
