// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: read.c.v
// Author: Fernando Martínez Santa - Stiven Cortazar Cortazar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: READ functions (Ai_Thinker_Ai-WB2-32S-Kit)
//              (PC port) 

module adc

#define adc__read(PIN_NAME)   analogRead(PIN_NAME)