// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: pin.c.v
// Author: Fernando Martínez Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: PIN functions (Ai_Thinker_Ai-WB2-32S-Kit)
//              (PC port) 

module pin

#define pin__out		OUTPUT
#define pin__in			INPUT
#define pin__in_pullup	INPUT_PULLUP

fn init() {

}