// Project Name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2022-2023
// License: MIT
//
// Description: Builtin definitions
//              (PC port) 
module main


enum Pin_names {    // enumerated type for the pin names
    gp0 = 0    
    gp1
    gp2
    gp3
    gp4
    gp5
    gp6
    gp7
    gp8
    gp9
    gp10
    gp11
    gp12
    gp13
    gp14
    gp15
    gp16
    gp17
    gp18
    gp19
    gp20
    gp21
    gp22
    gp23
    gp24
    gp25
    gp26
    gp27
    gp28
    gp29
}

enum Builtin_names {
	led0 = 25
}

enum Pin_modes {
	input = 0
	output
	in_pullup
}

enum ADC_pin_names {
	a0 = 14
	a1
	a2
	a3
	a4
	a5
	a6
	a7
}
