// Project Name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Pin-port functions
module port

// Port names
@[as_macro] pub const b = 0
@[as_macro] pub const c = 1
@[as_macro] pub const d = 2
// @[as_macro] pub const e = 3
// @[as_macro] pub const f = 4
// @[as_macro] pub const g = 5
// @[as_macro] pub const h = 6
// @[as_macro] pub const j = 7
// @[as_macro] pub const k = 8
// @[as_macro] pub const l = 9

@[as_macro] pub const all_inputs = 0b11111111
@[as_macro] pub const all_outputs = 0b00000000