module pic12f6xx

pub const description = 'API for the PIC12F6xx family devices'
