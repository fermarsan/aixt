module adc
fn init(){

}