// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: uart.c.v
// Author: Fernando Martínez Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: UART functions (Ai_Thinker_Ai-WB2-32S-Kit)
//              (PC port) 

<<<<<<< HEAD
fn init() {

}
=======
module uart
>>>>>>> eb738258f8b308832f65c20f9d5f8c2af4249322
