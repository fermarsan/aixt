module uart

#define uart__setup(BAUND_RATE)		Serial.begin(BAUND_RATE)
fn.init(){

}