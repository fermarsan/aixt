module time

#define time.sleep_ms(TIME)  delay(TIME)
