module uart

#define	uart__any()		RCIF