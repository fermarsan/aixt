// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git
// File Name: adc.c.v
// Author: Fernando Martinez Santa - Arley Junco - Luis Quevedo 
// Date: 2024
// License : MIT

module  adc

fn init() {
	
}