// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2023-2024
// License: MIT
//
// Description: input and printing functions.
module uart

#include <stdio.h>
#include <string.h>
	
fn C.init()