module uart

#define uart__ready()		Serial.available()