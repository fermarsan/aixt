// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git

// Author: Farith Ochoa León, Delipe Cardozo and Fernando M. Santa 
// License : MIT

module pwm 

#define pwm.write(PIN, VALUE) 			  analogWrite(PIN, VALUE)