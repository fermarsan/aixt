module xc16

pub const description = 'Workspace for the xc16 compiler modules'
