// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Pin management functions Arduino devices
module pin

// pin names
pub const d0   = 0    
pub const d1   = 1
pub const d2   = 2
pub const d3   = 3
pub const d4   = 4
pub const d5   = 5
pub const d6   = 6
pub const d7   = 7
pub const d8   = 8
pub const d9   = 9
pub const d10  = 10
pub const d11  = 11
pub const d12  = 12
pub const d13  = 13


// pin modes
pub const input		= 0
pub const output	= 1
pub const in_pullup = 2
