module main

#include "CH57x_common.h"
#define true 1

fn init() {
	//SetSysClock(CLK_SOURCE_PLL_60MHz)
}
