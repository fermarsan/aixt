// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2025
// License: MIT
//
// Description: Aixt's builtin components module
module builtin

// eprint adds a new error message to stderr (Aixt's table error list).
// This function does not generate any code
pub fn eprint(msg string)