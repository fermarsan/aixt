module uart
fn init(){

}