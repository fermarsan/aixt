module time
fn_init(){

}