// Author: Luis Alfredo Pinto Medina and Fernando M. Santa
// Date: 2024
//
// ## Description
// Builtin definitions (PIC16F88x port)

module main

#include <xc.h>
#include <stdio.h>
#include <stdbool.h>
#include <stdint.h>

#include "builtin.c"
