module pwm
fn.init(){

}