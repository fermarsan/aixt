// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: 
// Date: 
// License: MIT
//
// Description: 
module time

#include <libpic30.h>	//(PIC24, dsPIC33)
