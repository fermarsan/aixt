// Project Name : Aixt: http://github.com/fermansan/aixt.git
// Author: Fernando M. Santa
// License : MIT
// Date: 2025
//
// ## Description
// ADC functions for ESP32C3-CORE
module adc


pub const ch0 = 0
pub const ch1 = 1
pub const ch2 = 2
pub const ch3 = 3
pub const ch4 = 4
