module time

#define time__sleep_us(TIME)	delayMicroseconds(TIME)
fn.init(){

}