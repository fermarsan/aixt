// Project name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2025
// License: MIT
//
// Description: External interrupts management functions for 12F family
module ext

#include "ext.c"

@[as_macro] pub const rising  = 1
@[as_macro] pub const falling = 0