// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git
// File Name: adc.c.v
// Author: Farith Ochoa León, Delipe Cardozo and Fernando Martinez Santa 
// License : MIT

module pwm 

#define pwm__write(PIN, VALUE) 			  analogWrite(PIN, VALUE)