module time

#define time__sleep(S)    delay(S*1000)