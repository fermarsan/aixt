module time

#define time.sleep_ms(TIME)	mtimer_delay_ms(TIME)