// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fabián A. Rojas Acosta, Alberto Pinzón Valero and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: PWM functions (LQFP32 MiniEVB Nano - LGT8F328P port)
module pwm

fn init() { //  init function call setup or initialization code

}