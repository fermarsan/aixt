// _File:_ https://github.com/fermarsan/aixt/blob/main/
// Authors:
//	 - Julian Camilo Guzmán Zambrano
//	 - Juan Pablo Gonzalez Penagos
//	 - Fernando M. Santa
//
// _Date:_ 2022-2024
//
// // ## Description
// PIN functions (Blue Pill_STM32F103C)
//              (PC port)

module pin

@[as_macro] pub const rx = u8(C.PA9)
@[as_macro] pub const tx = u8(C.PA10)
@[as_macro] pub const p1 = u8(C.PA0)
@[as_macro] pub const p2 = u8(C.PA1)
@[as_macro] pub const p3 = u8(C.PA2)
@[as_macro] pub const p4 = u8(C.PA3)
@[as_macro] pub const p5 = u8(C.PA4)
@[as_macro] pub const p6 = u8(C.PA5)
@[as_macro] pub const p7 = u8(C.PA6)
@[as_macro] pub const p8 = u8(C.PA7)
@[as_macro] pub const p9 = u8(C.PA8)
@[as_macro] pub const p10 = u8(C.PA13)
@[as_macro] pub const p11 = u8(C.PA14)
@[as_macro] pub const p12 = u8(C.PA15)
@[as_macro] pub const p13 = u8(C.PB0)
@[as_macro] pub const p14 = u8(C.PB1)
@[as_macro] pub const p15 = u8(C.PB2)
@[as_macro] pub const p16 = u8(C.PB3)
@[as_macro] pub const p17 = u8(C.PB4)
@[as_macro] pub const p18 = u8(C.PB5)
@[as_macro] pub const p19 = u8(C.PB6)
@[as_macro] pub const p20 = u8(C.PB7)
@[as_macro] pub const p21 = u8(C.PB8)
@[as_macro] pub const p22 = u8(C.PB9)
@[as_macro] pub const p23 = u8(C.PB10)
@[as_macro] pub const p24 = u8(C.PB11)
@[as_macro] pub const p25 = u8(C.PB12)
@[as_macro] pub const p26 = u8(C.PB13)
@[as_macro] pub const p27 = u8(C.PB14)
@[as_macro] pub const p28 = u8(C.PB15)
