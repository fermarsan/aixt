module pin

#define pin__out		OUTPUT
#define pin__in			INPUT
#define pin__in_pullup	INPUT_PULLUP

fn init() {

}