// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: Pin port management functions (Explorer16-PIC24 port)
module port


fn init() {
	
}