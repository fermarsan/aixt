module PIC18

pub const description = 'Workspace for the PIC18 family devices'
