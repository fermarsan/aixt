// Project name: Aixt https://github.com/fermarsan/aixt.git
// Authors:
//	 - Julian Camilo Guzmán Zambrano
//	 - Juan Pablo Gonzalez Penagos
//	 - Fernando M. Santa
// Date: 2022-2025
// License: MIT
//
// Description: ADC functions
module adc

// adc channels
pub const ch0 = u8(C.PA0)
pub const ch1 = u8(C.PA1)
pub const ch2 = u8(C.PA2)
pub const ch3 = u8(C.PA3)
pub const ch4 = u8(C.PA4)
pub const ch5 = u8(C.PA5)
pub const ch6 = u8(C.PA6)
pub const ch7 = u8(C.PA7)
pub const ch8 = u8(C.PB0)
pub const ch9 = u8(C.PB1)