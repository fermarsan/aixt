// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: 
// Date: 
// License: MIT
module time

// sleep_us is a delay function in microseconds for the Aixt Explorer16-PIC24 port. 
#define time__sleep_us(TIME)    __delay_us(TIME)