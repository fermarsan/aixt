module pic16f87x

pub const description = 'API for the PIC16F87x family devices'
