// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: read_1.c.v
// Author: Fernando Martínez Santa - Julian Camilo Guzmán Zambrano - Juan Pablo Gonzalez Penagos
// Date: 2022-2024
// License: MIT
//
// // Description: READ_1 functions (Blue Pill_STM32F103C)
//              (PC port) 

module uart

#define uart__read_1   Serial1.read