// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024-2025
//
// ## Description
// Pin port management functions (Exp16-PIC24 port)
module port

@[as_macro] pub const a = 0 // port ids
@[as_macro] pub const b = 1
@[as_macro] pub const c = 2
@[as_macro] pub const d = 3
@[as_macro] pub const e = 4
@[as_macro] pub const f = 5
@[as_macro] pub const g = 6
