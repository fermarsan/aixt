module time

#define time.sleep(TIME) delay(TIME*1000)
