// ## Description
// This is a workspace for the Microchip devices
module PIC16_generic

pub const description = 'Workspace for the PIC16 family devices'
