// Author: Fernando M. Santa - Daniel Polo - Edwin Barrera - Javier Leon - Camilo Lucas
// Date: 2022-2025
//
// ## Description
// pwm write functions (CY8CKIT-049-42XX)

module pwm

// @[as_macro]
// pub fn write(channel any, val any) {
// 	C.PWM_WRITE(channel, val)
// }

@[as_macro]
pub fn write(channel int, val any) {
	match channel {
		pwm.ch0 {
			C.pwm0_WriteCompare(val)
		}
		pwm.ch1 {
			C.pwm1_WriteCompare(val)
		}
		pwm.ch2 {
			C.pwm2_WriteCompare(val)
		}
		else { }
	}
}
