// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Builtin definitions (Arduino Uno - ATmega328P port)
module main

#include "builtin.c"

@[as_macro]	const led_0 = 13
