module Arduino

pub const description = 'Arduino targets workspace'
