// Project name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2022-2025
// License: MIT
//
// Description: Builtin definitions (XIAO-SAM21 port) 
module main
