module uart
fn_init(){

}