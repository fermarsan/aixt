module adc
fn_init(){

}