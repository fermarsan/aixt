// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
//
// ## Description
// PWM functions (Exp16-PIC24 port)
module pwm



fn C.write(duty u8)
