module uart

#define uart__setup(BAUD_RATE)   Serial.begin(BAUD_RATE)