// Author: Fernando M. Santa
// Date: 2024

module lcd

// print function prints data to the serial port as human-readable ASCII text
@[as_macro]
pub fn setup(p1 u8,p2 u8) {
C.LCD_BEGIN(p1,p2)
}
