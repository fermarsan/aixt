// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: sleep_us.c.v
// Author: Fernando Martínez Santa - Stiven Cortazar Cortazar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: SLEEP_us functions (Ai_Thinker_Ai-WB2-32S-Kit)
//              (PC port) 

module time

#define time__sleep_us(US)    delayMicroseconds(US)