// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git

// Author: Farith Ochoa León, Delipe Cardozo and Fernando M. Santa 
// License : MIT

module adc 

#define adc.read(PIN_NAME) 	 	analogRead(PIN_NAME)
