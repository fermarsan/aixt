// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: outpwm.c.v
// Author: Fernando M. Santa - Johann Escobar Guzmán - Daniel Andrés Vásquez Gómez
// Date: 2023-2024
// License: MIT
//
// // Description: out functions (W801)
//              (PC port) 

module pin

#define PWM__OUT  PWM_OUT