// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: uart.c.v
// Author: Fernando M. Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: fn init() functions (Ai_Thinker_Ai-WB2-32S-Kit)

module uart

fn init() {

}