module exp16_pic24

pub const description = 'API for the Exp16_PIC24 family devices'
