// Author: Fernando M. Santa
// Date: 2022-2023
//
// ## Description
// Builtin definitions
//              (PC port)
module main

// builtin LED
const led0 = 25
