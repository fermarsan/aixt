// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: pwm.c.v
// Author: Fernando Martínez Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// // Description: PWM functions (Ai_Thinker_Ai-WB2-32S-Kit)
//              (PC port) 

module pwm

fn init() {

}