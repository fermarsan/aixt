module time
fn init() {

}
