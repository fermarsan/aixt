module PIC16

pub const description = 'Workspace for the PIC16 family devices'
