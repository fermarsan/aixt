<<<<<<< HEAD
// Project name: Aixt https://github.com/fermarsan/aixt.git
// Authors:
//	 - Julian Camilo Guzmán Zambrano
//	 - Juan Pablo Gonzalez Penagos
//	 - Fernando M. Santa
// Date: 2022-2024
// License: MIT
//
// // Description: ADC functions (Blue Pill_STM32F103C)
//              (PC port) 

module adc
=======
module adc


>>>>>>> d4993b91b137dd499e1bd8c91cce3c82d74f8e77
