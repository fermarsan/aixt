// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: builtin.c.v
// Author: Fernando M. Santa - Johann Escobar Guzmán - Daniel Andrés Vásquez Gómez
// Date: 2023-2024
// License: MIT
//
// Description: Builtin definitions
//              (PC port) 
module main

enum __pin_names {    // enumerated type for the pin names

led1 = LED_BUILTIN_1
led2 = LED_BUILTIN_2
led3 = LED_BUILTIN_3
led4 = LED_BUILTIN_4
led5 = LED_BUILTIN_5
led6 = LED_BUILTIN_6
led7 = LED_BUILTIN_7

a1 = PB21
a2 = PB22
a3 = PB23
a4 = PB24
a5 = PB0
a6 = PB1



pin1 = PB21
pin2 = PB22

}

fn init() {

}
