// Project Name : Aixt: http://github.com/fermansan/aixt.git
// Authors:
//	- Farith Ochoa Leon
//	- Felipe Cardozo
//	- Fernando M. Santa
// Date: 2024
// License : MIT

module uart 

