module api

pub const description = 'API workspace for PIC16F87x'
