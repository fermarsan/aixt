// Author: Fernando M. Santa
// Date: 29/01/2025
//
// ## Description
// Example of a Library module.
//
module ex_array

fn C.ArrayMin(src []any, idx u16, len u16) any
