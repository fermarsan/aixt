// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2023-2024
// License: MIT
module cgen2

// init_output_file initializes the output file stream.
fn (mut gen Gen) init_output_file() {
	mut c_line := ''
	c_line += '// This '
    c_line += match gen.setup.backend {
		'nxc' 		{ 'NXC ' }
		'arduino'	{ 'Arduino ' }  
		else 		{ 'C ' }
	}
    gen.out << c_line + 'code was automatically generated by Aixt Project'
	gen.out << '//     https://github.com/fermarsan/aixt'
	gen.out << '// Device = ${gen.setup.device}'
	gen.out << '// Board = ${gen.setup.board}'
	gen.out << '// Backend = ${gen.setup.backend}\n'

	gen.out << '\n___preprocessor_block___' 

	for v_type, c_type in gen.setup.compiler_types {	// type definitions
		// println('>>>>>>>>>>>>>>>>>> ${c_type} , ${v_type}==================')
		if c_type != v_type {
			gen.out << if v_type == 'int' {
				'typedef ${c_type} i32;'
			} else if c_type == 'NOT SUPPORTED' {
				'// typedef ${c_type} ${v_type};'
			} else if gen.setup.backend == 'arduino' && v_type == "u16" {
				'// typedef ${c_type} ${v_type};'
			} else {
				'typedef ${c_type} ${v_type};'
			}
		}
	} 
	// gen.out += '\n___includes_block___\n'
	// gen.out += '\n___macros_block___\n' 
	gen.out << '\n___definitions_block___\n'
}