// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Cristian Garzón
// Date: 2023 - 2024
// Description: UART functions (WCH-CH573F)

module uart

@[inline]
pub fn uart.write(DATA) {
	C.R8_UART0_THR = DATA
}