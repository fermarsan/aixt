// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: builtin.c
// Author: Fernando Martínez Santa - Julian Camilo Guzmán Zambrano - Juan Pablo Gonzalez Penagos
// Date: 2022-2023
// License: MIT
//
// Description: Builtin definitions
//              (PC port) 
module main

enum __pin_names {    // enumerated type for the pin names
 
    RX=PA11
    TX=PA10
    PA0
    PA1
    PA2
    PA3
    PA4
    PA5
    PA6
    PA7
    PB0
    PB1
    PB10
    PB11
    PB12
    PB13
    PB14
    PB15
    PA8
    PB3
    PB4
    PB5
    PB6
    PB7
    PB8
    PB9

}

fn init() {

}
