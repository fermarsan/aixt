// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2025
// License: MIT
//
// Description: lcd module (Arduino Nano - ATmega328P port)
module disp7seg

#include "disp7seg.c"


fn C.DISP7SEG_BEGIN() void
fn C.DISP7SEG_SETVALUE(P1 int) 
fn C.DISP7SEG_SETPRECISION(P1 int) 
fn C.DISP7SEG_SETLEADINGZEROS(P1 bool) 
fn C.DISP7SEG_SETBLANK(P1 bool) 
fn C.DISP7SEG_SETDIGIT(P1 int, P2 int) 
fn C.DISP7SEG_SETDECIMALPOINT(P1 int, P2 bool) 





