// Project Name: Aixt project https://gitlab.com/fermarsan/aixt-project.git
// File Name: builtin.c.v
// Author: Fernando Martínez Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2023
// License: MIT
//
// Description: Builtin definitions

module main

enum __pin_names {    // enumerated type for the pin names
    IO11=11
    IO14=14
    IO17=17
    IO3=3
    IO4=4
    IO5=5
    RX=7
    TX=16
    IO12=12

}

fn init() {

}
