// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// File Name: uart.c.v
// Author: Jan Carlo Peñuela Jurado and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: uart
//              (PIC18F452)
module uart

#include <xc.h>

fn init() {
    
}