module my_sub

// add (integer)
pub fn add(x int, y int) int {
	return x + y
}