// Project Nme : Aixt project : http://gitlab.com/fermansan/aixt-project.git
// File Name: adc.c.v
// Author: Farith Ochoa León, Delipe Cardozo and Fernando M. Santa 
// License : MIT

module pin 

#define pin__output 		OUTPUT 
#define pin__input 			INPUT
#define pin__input_pullup 	INPUT_PULLUP

fn init () { 
	
}