module uart

#define uart__available(MESSAGE)	Serial.available(MESSAGE)