// Project Name : Aixt: http://github.com/fermansan/aixt.git
//
// _Author:_ Farith Ochoa León, Delipe Cardozo and Fernando M. Santa 
// License : MIT
//
// _Date:_ 2024-2025
//
// ## Description
// ADC functions
module adc

// ADC pin names
pub const ch0 = 0
pub const ch1 = 1
pub const ch2 = 2
pub const ch3 = 3
pub const ch4 = 4