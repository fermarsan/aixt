// Project Name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa - Julian Camilo Guzmán Zambrano - Juan Pablo Gonzalez Penagos
// Date: 2022-2024
// License: MIT
//
// // Description: PIN functions (Blue Pill_STM32F103C)
//              (PC port) 

module pin

#define output		OUTPUT
#define input		INPUT
#define in_pullup	INPUT_PULLUP

fn init() {

}