module uart

#define uart__read_1()		Serial1.read()
