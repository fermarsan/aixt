// Author: Cristian Garzón
// Date: 2023 - 2024
// ## Description
// UART1 functions (WCH-CH573F)

module uart1

fn C.print(msg string)