module time

#define time.sleep(S)    delay(S*1000)