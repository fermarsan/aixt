// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Andrés Felipe Fajardo Duarte and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: UART management functions  (PIC18F2550 port)

module uart

fn read() rune{
  return RCREG
}