module time

#define time__sleep(TIME) delay(TIME*1000)
fn.init(){

}