module time

#define time.sleep(TIME) delay(TIME*1000)

#define time.sleep_ms(TIME)  delay(TIME)

#define time.sleep_us(TIME)	delayMicroseconds(TIME)