module adc

#define adc__read(PIN_NAME)   analogRead(PIN_NAME)