// Project Name: Aixt, https://github.com/fermarsan/aixt.git

// Author: Jan Carlo Peñuela Jurado and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: Pin management functions (PIC18F452)
module pin

#include <xc.h>

#define output 0   // pin mode (direction)
#define input  1

fn init() {
    
}