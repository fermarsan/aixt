module main


fn init() {
	
}