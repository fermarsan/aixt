// Project name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa - Stiven Cortázar Cortázar - Yesid Reyes Tique
// Date: 2022-2024
// License: MIT
//
// Description: pin functions (Ai_Thinker_Ai-WB2-32S-Kit)

module pin

//  pin names
pub const gpio11 = 11
pub const gpio14 = 14
pub const gpio17 = 17
pub const gpio3  = 3
pub const gpio4  = 4
pub const gpio5  = 5
pub const gpio7  = 7
pub const gpio16 = 16
pub const gpio12 = 12

