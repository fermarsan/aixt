// Project name: Aixt, https://github.com/fermarsan/aixt.git
//
// _Author:_ Fernando M. Santa
//
// _Date:_ 29/01/2025
//
// ## Description
// Example of a Library module.
//
module ex_array

