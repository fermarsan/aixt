// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// File Name: time.c.v
// Author: Andrés Felipe Fajardo Duarte and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: TIME delay function
//              (PIC18F2550)

module time

#include <xc.h>

fn init() {
    
}