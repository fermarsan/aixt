// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024-2025
// License: MIT
//
// Description: Pin management functions Arduino devices
module pin_fn

// pin names 
@[as_macro] pub const d0 = 0 
@[as_macro] pub const d1 = 1
@[as_macro] pub const d2 = 2
@[as_macro] pub const d3 = 3
@[as_macro] pub const d4 = 4
@[as_macro] pub const d5 = 5
@[as_macro] pub const d6 = 6
@[as_macro] pub const d7 = 7
@[as_macro] pub const d8 = 8
@[as_macro] pub const d9 = 9
@[as_macro] pub const d10 = 10
@[as_macro] pub const d11 = 11
@[as_macro] pub const d12 = 12
@[as_macro] pub const d13 = 13
@[as_macro] pub const d14 = 14
@[as_macro] pub const d15 = 15
@[as_macro] pub const d16 = 16
@[as_macro] pub const d17 = 17
@[as_macro] pub const d18 = 18
@[as_macro] pub const d19 = 19
@[as_macro] pub const d22 = 22 
@[as_macro] pub const d23 = 23
@[as_macro] pub const d24 = 24
@[as_macro] pub const d25 = 25
@[as_macro] pub const d26 = 26
@[as_macro] pub const d27 = 27
@[as_macro] pub const d28 = 28
@[as_macro] pub const d29 = 29
@[as_macro] pub const d30 = 30
@[as_macro] pub const d31 = 31
@[as_macro] pub const d32 = 32
@[as_macro] pub const d33 = 33
@[as_macro] pub const d34 = 34
@[as_macro] pub const d35 = 35
@[as_macro] pub const d36 = 36
@[as_macro] pub const d37 = 37
@[as_macro] pub const d38 = 38
@[as_macro] pub const d39 = 39
@[as_macro] pub const d40 = 40
@[as_macro] pub const d41 = 41
@[as_macro] pub const d42 = 42
@[as_macro] pub const d43 = 43
@[as_macro] pub const d44 = 44
@[as_macro] pub const d45 = 45
@[as_macro] pub const d46 = 46
@[as_macro] pub const d47 = 47
@[as_macro] pub const d48 = 48
@[as_macro] pub const d49 = 49
@[as_macro] pub const d50 = 50
@[as_macro] pub const d51 = 51
@[as_macro] pub const d52 = 52
@[as_macro] pub const d53 = 53
@[as_macro] pub const d54 = 54
@[as_macro] pub const d55 = 55
@[as_macro] pub const d56 = 56
@[as_macro] pub const d57 = 57
@[as_macro] pub const d58 = 58
@[as_macro] pub const d59 = 59
@[as_macro] pub const d60 = 60
@[as_macro] pub const d61 = 61
@[as_macro] pub const d62 = 62
@[as_macro] pub const d63 = 63
@[as_macro] pub const d64 = 64
@[as_macro] pub const d65 = 65
@[as_macro] pub const d66 = 66
@[as_macro] pub const d67 = 67
@[as_macro] pub const d68 = 68
@[as_macro] pub const d69 = 69


// builtin LED
@[as_macro]	pub const led0 = 13

fn init() {
	setup(led0, pin_fn.output)
}