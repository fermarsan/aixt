// Project name: Aixt project, https://github.com/fermarsan/aixt.git
// Authors: Fernando M. Santa
// Date: 2025
// License: MIT
//
// Description: Builtin definitions PIC12F6xx

module main

#include <xc.h>
#include <stdint.h>
#include <stdbool.h>

#include "builtin.c"
