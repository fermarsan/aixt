// Project Name: Aixt project, https://github.com/fermarsan/aixt.git
// Author: Luis Alfredo Pinto Medina and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: Pin-port functions (PIC16F886 port)

module port

#define TRISa	TRISA	// port setup name equivalents
#define TRISb	TRISB
#define TRISc	TRISC

#define PORTa	PORTA	// port in name equivalents
#define PORTb	PORTB
#define PORTc	PORTC

#define	port__all_inputs	0xFF	// port mode constants
#define	port__all_outputs	0x00

