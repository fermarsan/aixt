// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fabián A. Rojas Acosta, Alberto Pinzón Valero and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: ADC functions (Arduino Nano - ATmega328P port)
module adc

pub const (
	a0 = 14
	a1 = 15
	a2 = 16
	a3 = 17
	a4 = 18
	a5 = 19
	a6 = 20
	a7 = 21
)