// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fabián A. Rojas Acosta, Alberto Pinzón Valero and Fernando Martínez Santa
// Date: 2024
// License: MIT
//
// Description: Pin management functions (Arduino Nano - ATmega328P port)
module pin

pub const (
	input = 0x0
	output = 0x1
	in_pullup = 0x2
)