// Project name: Aixt, https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa
// Date: 2024
//
// ## Description
// Pin management Nucleo-L031K6
module pin

// pin names
@[as_macro] pub const d0   = 0    
@[as_macro] pub const d1   = 1
@[as_macro] pub const d2   = 2
@[as_macro] pub const d3   = 3
@[as_macro] pub const d4   = 4
@[as_macro] pub const d5   = 5
@[as_macro] pub const d6   = 6
@[as_macro] pub const d7   = 7
@[as_macro] pub const d8   = 8
@[as_macro] pub const d9   = 9
@[as_macro] pub const d10  = 10
@[as_macro] pub const d11  = 11
@[as_macro] pub const d12  = 12
@[as_macro] pub const d13  = 13
