// module importing

import time { sleep }
import machine

mut a := 0.0

for {
	sleep(1)
	a++
}