// Project Name: Aixt https://github.com/fermarsan/aixt.git
// Author: Fernando M. Santa - Daniel Polo - Edwin Barrera - Javier Leon - Camilo Lucas
// Date: 2022-2025
// License: MIT
//
// // Description: adc functions (CY8CKIT-049-42XX)

module adc

fn C.adc_Start()
fn C.adc_StartConvert()




