module sw_uart

#define sw_uart.setup(BAUDRATE)	sw_uart.baudrate = BAUDRATE