// Project Name: Aixt, https://github.com/fermarsan/aixt.git
// File Name: adc.c.v
// Author: Andrés Felipe Fajardo Duarte and Fernando M. Santa
// Date: 2024
// License: MIT
//
// Description: ADC management functions  (PIC18F2550 port)

module adc

#include <xc.h>

fn init() {
    
}